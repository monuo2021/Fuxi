module GHR(
  input        clock,
  input        io_branch,
  input        io_taken,
  output [4:0] io_ghr
);
  reg [4:0] ghr; // @[GHR.scala 23:16]
  reg [31:0] _RAND_0;
  wire [4:0] _T_1 = {ghr[3:0],io_taken}; // @[Cat.scala 30:58]
  assign io_ghr = ghr; // @[GHR.scala 29:10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ghr = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (io_branch) begin
      ghr <= _T_1;
    end
  end
endmodule
module PHT(
  input        clock,
  input        reset,
  input        io_lastBranch,
  input        io_lastTaken,
  input  [4:0] io_lastIndex,
  input  [4:0] io_index,
  output       io_taken
);
  reg [1:0] counters_0; // @[PHT.scala 23:26]
  reg [31:0] _RAND_0;
  reg [1:0] counters_1; // @[PHT.scala 23:26]
  reg [31:0] _RAND_1;
  reg [1:0] counters_2; // @[PHT.scala 23:26]
  reg [31:0] _RAND_2;
  reg [1:0] counters_3; // @[PHT.scala 23:26]
  reg [31:0] _RAND_3;
  reg [1:0] counters_4; // @[PHT.scala 23:26]
  reg [31:0] _RAND_4;
  reg [1:0] counters_5; // @[PHT.scala 23:26]
  reg [31:0] _RAND_5;
  reg [1:0] counters_6; // @[PHT.scala 23:26]
  reg [31:0] _RAND_6;
  reg [1:0] counters_7; // @[PHT.scala 23:26]
  reg [31:0] _RAND_7;
  reg [1:0] counters_8; // @[PHT.scala 23:26]
  reg [31:0] _RAND_8;
  reg [1:0] counters_9; // @[PHT.scala 23:26]
  reg [31:0] _RAND_9;
  reg [1:0] counters_10; // @[PHT.scala 23:26]
  reg [31:0] _RAND_10;
  reg [1:0] counters_11; // @[PHT.scala 23:26]
  reg [31:0] _RAND_11;
  reg [1:0] counters_12; // @[PHT.scala 23:26]
  reg [31:0] _RAND_12;
  reg [1:0] counters_13; // @[PHT.scala 23:26]
  reg [31:0] _RAND_13;
  reg [1:0] counters_14; // @[PHT.scala 23:26]
  reg [31:0] _RAND_14;
  reg [1:0] counters_15; // @[PHT.scala 23:26]
  reg [31:0] _RAND_15;
  reg [1:0] counters_16; // @[PHT.scala 23:26]
  reg [31:0] _RAND_16;
  reg [1:0] counters_17; // @[PHT.scala 23:26]
  reg [31:0] _RAND_17;
  reg [1:0] counters_18; // @[PHT.scala 23:26]
  reg [31:0] _RAND_18;
  reg [1:0] counters_19; // @[PHT.scala 23:26]
  reg [31:0] _RAND_19;
  reg [1:0] counters_20; // @[PHT.scala 23:26]
  reg [31:0] _RAND_20;
  reg [1:0] counters_21; // @[PHT.scala 23:26]
  reg [31:0] _RAND_21;
  reg [1:0] counters_22; // @[PHT.scala 23:26]
  reg [31:0] _RAND_22;
  reg [1:0] counters_23; // @[PHT.scala 23:26]
  reg [31:0] _RAND_23;
  reg [1:0] counters_24; // @[PHT.scala 23:26]
  reg [31:0] _RAND_24;
  reg [1:0] counters_25; // @[PHT.scala 23:26]
  reg [31:0] _RAND_25;
  reg [1:0] counters_26; // @[PHT.scala 23:26]
  reg [31:0] _RAND_26;
  reg [1:0] counters_27; // @[PHT.scala 23:26]
  reg [31:0] _RAND_27;
  reg [1:0] counters_28; // @[PHT.scala 23:26]
  reg [31:0] _RAND_28;
  reg [1:0] counters_29; // @[PHT.scala 23:26]
  reg [31:0] _RAND_29;
  reg [1:0] counters_30; // @[PHT.scala 23:26]
  reg [31:0] _RAND_30;
  reg [1:0] counters_31; // @[PHT.scala 23:26]
  reg [31:0] _RAND_31;
  wire [1:0] _GEN_1 = 5'h1 == io_lastIndex ? counters_1 : counters_0; // @[PHT.scala 27:34]
  wire [1:0] _GEN_2 = 5'h2 == io_lastIndex ? counters_2 : _GEN_1; // @[PHT.scala 27:34]
  wire [1:0] _GEN_3 = 5'h3 == io_lastIndex ? counters_3 : _GEN_2; // @[PHT.scala 27:34]
  wire [1:0] _GEN_4 = 5'h4 == io_lastIndex ? counters_4 : _GEN_3; // @[PHT.scala 27:34]
  wire [1:0] _GEN_5 = 5'h5 == io_lastIndex ? counters_5 : _GEN_4; // @[PHT.scala 27:34]
  wire [1:0] _GEN_6 = 5'h6 == io_lastIndex ? counters_6 : _GEN_5; // @[PHT.scala 27:34]
  wire [1:0] _GEN_7 = 5'h7 == io_lastIndex ? counters_7 : _GEN_6; // @[PHT.scala 27:34]
  wire [1:0] _GEN_8 = 5'h8 == io_lastIndex ? counters_8 : _GEN_7; // @[PHT.scala 27:34]
  wire [1:0] _GEN_9 = 5'h9 == io_lastIndex ? counters_9 : _GEN_8; // @[PHT.scala 27:34]
  wire [1:0] _GEN_10 = 5'ha == io_lastIndex ? counters_10 : _GEN_9; // @[PHT.scala 27:34]
  wire [1:0] _GEN_11 = 5'hb == io_lastIndex ? counters_11 : _GEN_10; // @[PHT.scala 27:34]
  wire [1:0] _GEN_12 = 5'hc == io_lastIndex ? counters_12 : _GEN_11; // @[PHT.scala 27:34]
  wire [1:0] _GEN_13 = 5'hd == io_lastIndex ? counters_13 : _GEN_12; // @[PHT.scala 27:34]
  wire [1:0] _GEN_14 = 5'he == io_lastIndex ? counters_14 : _GEN_13; // @[PHT.scala 27:34]
  wire [1:0] _GEN_15 = 5'hf == io_lastIndex ? counters_15 : _GEN_14; // @[PHT.scala 27:34]
  wire [1:0] _GEN_16 = 5'h10 == io_lastIndex ? counters_16 : _GEN_15; // @[PHT.scala 27:34]
  wire [1:0] _GEN_17 = 5'h11 == io_lastIndex ? counters_17 : _GEN_16; // @[PHT.scala 27:34]
  wire [1:0] _GEN_18 = 5'h12 == io_lastIndex ? counters_18 : _GEN_17; // @[PHT.scala 27:34]
  wire [1:0] _GEN_19 = 5'h13 == io_lastIndex ? counters_19 : _GEN_18; // @[PHT.scala 27:34]
  wire [1:0] _GEN_20 = 5'h14 == io_lastIndex ? counters_20 : _GEN_19; // @[PHT.scala 27:34]
  wire [1:0] _GEN_21 = 5'h15 == io_lastIndex ? counters_21 : _GEN_20; // @[PHT.scala 27:34]
  wire [1:0] _GEN_22 = 5'h16 == io_lastIndex ? counters_22 : _GEN_21; // @[PHT.scala 27:34]
  wire [1:0] _GEN_23 = 5'h17 == io_lastIndex ? counters_23 : _GEN_22; // @[PHT.scala 27:34]
  wire [1:0] _GEN_24 = 5'h18 == io_lastIndex ? counters_24 : _GEN_23; // @[PHT.scala 27:34]
  wire [1:0] _GEN_25 = 5'h19 == io_lastIndex ? counters_25 : _GEN_24; // @[PHT.scala 27:34]
  wire [1:0] _GEN_26 = 5'h1a == io_lastIndex ? counters_26 : _GEN_25; // @[PHT.scala 27:34]
  wire [1:0] _GEN_27 = 5'h1b == io_lastIndex ? counters_27 : _GEN_26; // @[PHT.scala 27:34]
  wire [1:0] _GEN_28 = 5'h1c == io_lastIndex ? counters_28 : _GEN_27; // @[PHT.scala 27:34]
  wire [1:0] _GEN_29 = 5'h1d == io_lastIndex ? counters_29 : _GEN_28; // @[PHT.scala 27:34]
  wire [1:0] _GEN_30 = 5'h1e == io_lastIndex ? counters_30 : _GEN_29; // @[PHT.scala 27:34]
  wire [1:0] _GEN_31 = 5'h1f == io_lastIndex ? counters_31 : _GEN_30; // @[PHT.scala 27:34]
  wire  _T_1 = _GEN_31 == 2'h3; // @[PHT.scala 27:34]
  wire  _T_2 = ~io_lastTaken; // @[PHT.scala 28:13]
  wire [1:0] _T_4 = _GEN_31 - 2'h1; // @[PHT.scala 29:58]
  wire  _T_5 = _GEN_31 == 2'h0; // @[PHT.scala 31:41]
  wire [1:0] _T_7 = _GEN_31 + 2'h1; // @[PHT.scala 33:58]
  wire [1:0] _GEN_353 = 5'h1 == io_index ? counters_1 : counters_0; // @[PHT.scala 46:33]
  wire [1:0] _GEN_354 = 5'h2 == io_index ? counters_2 : _GEN_353; // @[PHT.scala 46:33]
  wire [1:0] _GEN_355 = 5'h3 == io_index ? counters_3 : _GEN_354; // @[PHT.scala 46:33]
  wire [1:0] _GEN_356 = 5'h4 == io_index ? counters_4 : _GEN_355; // @[PHT.scala 46:33]
  wire [1:0] _GEN_357 = 5'h5 == io_index ? counters_5 : _GEN_356; // @[PHT.scala 46:33]
  wire [1:0] _GEN_358 = 5'h6 == io_index ? counters_6 : _GEN_357; // @[PHT.scala 46:33]
  wire [1:0] _GEN_359 = 5'h7 == io_index ? counters_7 : _GEN_358; // @[PHT.scala 46:33]
  wire [1:0] _GEN_360 = 5'h8 == io_index ? counters_8 : _GEN_359; // @[PHT.scala 46:33]
  wire [1:0] _GEN_361 = 5'h9 == io_index ? counters_9 : _GEN_360; // @[PHT.scala 46:33]
  wire [1:0] _GEN_362 = 5'ha == io_index ? counters_10 : _GEN_361; // @[PHT.scala 46:33]
  wire [1:0] _GEN_363 = 5'hb == io_index ? counters_11 : _GEN_362; // @[PHT.scala 46:33]
  wire [1:0] _GEN_364 = 5'hc == io_index ? counters_12 : _GEN_363; // @[PHT.scala 46:33]
  wire [1:0] _GEN_365 = 5'hd == io_index ? counters_13 : _GEN_364; // @[PHT.scala 46:33]
  wire [1:0] _GEN_366 = 5'he == io_index ? counters_14 : _GEN_365; // @[PHT.scala 46:33]
  wire [1:0] _GEN_367 = 5'hf == io_index ? counters_15 : _GEN_366; // @[PHT.scala 46:33]
  wire [1:0] _GEN_368 = 5'h10 == io_index ? counters_16 : _GEN_367; // @[PHT.scala 46:33]
  wire [1:0] _GEN_369 = 5'h11 == io_index ? counters_17 : _GEN_368; // @[PHT.scala 46:33]
  wire [1:0] _GEN_370 = 5'h12 == io_index ? counters_18 : _GEN_369; // @[PHT.scala 46:33]
  wire [1:0] _GEN_371 = 5'h13 == io_index ? counters_19 : _GEN_370; // @[PHT.scala 46:33]
  wire [1:0] _GEN_372 = 5'h14 == io_index ? counters_20 : _GEN_371; // @[PHT.scala 46:33]
  wire [1:0] _GEN_373 = 5'h15 == io_index ? counters_21 : _GEN_372; // @[PHT.scala 46:33]
  wire [1:0] _GEN_374 = 5'h16 == io_index ? counters_22 : _GEN_373; // @[PHT.scala 46:33]
  wire [1:0] _GEN_375 = 5'h17 == io_index ? counters_23 : _GEN_374; // @[PHT.scala 46:33]
  wire [1:0] _GEN_376 = 5'h18 == io_index ? counters_24 : _GEN_375; // @[PHT.scala 46:33]
  wire [1:0] _GEN_377 = 5'h19 == io_index ? counters_25 : _GEN_376; // @[PHT.scala 46:33]
  wire [1:0] _GEN_378 = 5'h1a == io_index ? counters_26 : _GEN_377; // @[PHT.scala 46:33]
  wire [1:0] _GEN_379 = 5'h1b == io_index ? counters_27 : _GEN_378; // @[PHT.scala 46:33]
  wire [1:0] _GEN_380 = 5'h1c == io_index ? counters_28 : _GEN_379; // @[PHT.scala 46:33]
  wire [1:0] _GEN_381 = 5'h1d == io_index ? counters_29 : _GEN_380; // @[PHT.scala 46:33]
  wire [1:0] _GEN_382 = 5'h1e == io_index ? counters_30 : _GEN_381; // @[PHT.scala 46:33]
  wire [1:0] _GEN_383 = 5'h1f == io_index ? counters_31 : _GEN_382; // @[PHT.scala 46:33]
  assign io_taken = _GEN_383[1]; // @[PHT.scala 46:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  counters_0 = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  counters_1 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  counters_2 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  counters_3 = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  counters_4 = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  counters_5 = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  counters_6 = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  counters_7 = _RAND_7[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  counters_8 = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  counters_9 = _RAND_9[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  counters_10 = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  counters_11 = _RAND_11[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  counters_12 = _RAND_12[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  counters_13 = _RAND_13[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  counters_14 = _RAND_14[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  counters_15 = _RAND_15[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  counters_16 = _RAND_16[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  counters_17 = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  counters_18 = _RAND_18[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  counters_19 = _RAND_19[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  counters_20 = _RAND_20[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  counters_21 = _RAND_21[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  counters_22 = _RAND_22[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  counters_23 = _RAND_23[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  counters_24 = _RAND_24[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  counters_25 = _RAND_25[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  counters_26 = _RAND_26[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  counters_27 = _RAND_27[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  counters_28 = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  counters_29 = _RAND_29[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  counters_30 = _RAND_30[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  counters_31 = _RAND_31[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      counters_0 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h0 == io_lastIndex) begin
            counters_0 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h0 == io_lastIndex) begin
            counters_0 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h0 == io_lastIndex) begin
          counters_0 <= _T_4;
        end
      end else if (5'h0 == io_lastIndex) begin
        counters_0 <= _T_7;
      end
    end
    if (reset) begin
      counters_1 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h1 == io_lastIndex) begin
            counters_1 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h1 == io_lastIndex) begin
            counters_1 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h1 == io_lastIndex) begin
          counters_1 <= _T_4;
        end
      end else if (5'h1 == io_lastIndex) begin
        counters_1 <= _T_7;
      end
    end
    if (reset) begin
      counters_2 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h2 == io_lastIndex) begin
            counters_2 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h2 == io_lastIndex) begin
            counters_2 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h2 == io_lastIndex) begin
          counters_2 <= _T_4;
        end
      end else if (5'h2 == io_lastIndex) begin
        counters_2 <= _T_7;
      end
    end
    if (reset) begin
      counters_3 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h3 == io_lastIndex) begin
            counters_3 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h3 == io_lastIndex) begin
            counters_3 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h3 == io_lastIndex) begin
          counters_3 <= _T_4;
        end
      end else if (5'h3 == io_lastIndex) begin
        counters_3 <= _T_7;
      end
    end
    if (reset) begin
      counters_4 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h4 == io_lastIndex) begin
            counters_4 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h4 == io_lastIndex) begin
            counters_4 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h4 == io_lastIndex) begin
          counters_4 <= _T_4;
        end
      end else if (5'h4 == io_lastIndex) begin
        counters_4 <= _T_7;
      end
    end
    if (reset) begin
      counters_5 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h5 == io_lastIndex) begin
            counters_5 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h5 == io_lastIndex) begin
            counters_5 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h5 == io_lastIndex) begin
          counters_5 <= _T_4;
        end
      end else if (5'h5 == io_lastIndex) begin
        counters_5 <= _T_7;
      end
    end
    if (reset) begin
      counters_6 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h6 == io_lastIndex) begin
            counters_6 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h6 == io_lastIndex) begin
            counters_6 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h6 == io_lastIndex) begin
          counters_6 <= _T_4;
        end
      end else if (5'h6 == io_lastIndex) begin
        counters_6 <= _T_7;
      end
    end
    if (reset) begin
      counters_7 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h7 == io_lastIndex) begin
            counters_7 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h7 == io_lastIndex) begin
            counters_7 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h7 == io_lastIndex) begin
          counters_7 <= _T_4;
        end
      end else if (5'h7 == io_lastIndex) begin
        counters_7 <= _T_7;
      end
    end
    if (reset) begin
      counters_8 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h8 == io_lastIndex) begin
            counters_8 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h8 == io_lastIndex) begin
            counters_8 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h8 == io_lastIndex) begin
          counters_8 <= _T_4;
        end
      end else if (5'h8 == io_lastIndex) begin
        counters_8 <= _T_7;
      end
    end
    if (reset) begin
      counters_9 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h9 == io_lastIndex) begin
            counters_9 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h9 == io_lastIndex) begin
            counters_9 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h9 == io_lastIndex) begin
          counters_9 <= _T_4;
        end
      end else if (5'h9 == io_lastIndex) begin
        counters_9 <= _T_7;
      end
    end
    if (reset) begin
      counters_10 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'ha == io_lastIndex) begin
            counters_10 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'ha == io_lastIndex) begin
            counters_10 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'ha == io_lastIndex) begin
          counters_10 <= _T_4;
        end
      end else if (5'ha == io_lastIndex) begin
        counters_10 <= _T_7;
      end
    end
    if (reset) begin
      counters_11 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'hb == io_lastIndex) begin
            counters_11 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'hb == io_lastIndex) begin
            counters_11 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'hb == io_lastIndex) begin
          counters_11 <= _T_4;
        end
      end else if (5'hb == io_lastIndex) begin
        counters_11 <= _T_7;
      end
    end
    if (reset) begin
      counters_12 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'hc == io_lastIndex) begin
            counters_12 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'hc == io_lastIndex) begin
            counters_12 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'hc == io_lastIndex) begin
          counters_12 <= _T_4;
        end
      end else if (5'hc == io_lastIndex) begin
        counters_12 <= _T_7;
      end
    end
    if (reset) begin
      counters_13 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'hd == io_lastIndex) begin
            counters_13 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'hd == io_lastIndex) begin
            counters_13 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'hd == io_lastIndex) begin
          counters_13 <= _T_4;
        end
      end else if (5'hd == io_lastIndex) begin
        counters_13 <= _T_7;
      end
    end
    if (reset) begin
      counters_14 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'he == io_lastIndex) begin
            counters_14 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'he == io_lastIndex) begin
            counters_14 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'he == io_lastIndex) begin
          counters_14 <= _T_4;
        end
      end else if (5'he == io_lastIndex) begin
        counters_14 <= _T_7;
      end
    end
    if (reset) begin
      counters_15 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'hf == io_lastIndex) begin
            counters_15 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'hf == io_lastIndex) begin
            counters_15 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'hf == io_lastIndex) begin
          counters_15 <= _T_4;
        end
      end else if (5'hf == io_lastIndex) begin
        counters_15 <= _T_7;
      end
    end
    if (reset) begin
      counters_16 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h10 == io_lastIndex) begin
            counters_16 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h10 == io_lastIndex) begin
            counters_16 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h10 == io_lastIndex) begin
          counters_16 <= _T_4;
        end
      end else if (5'h10 == io_lastIndex) begin
        counters_16 <= _T_7;
      end
    end
    if (reset) begin
      counters_17 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h11 == io_lastIndex) begin
            counters_17 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h11 == io_lastIndex) begin
            counters_17 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h11 == io_lastIndex) begin
          counters_17 <= _T_4;
        end
      end else if (5'h11 == io_lastIndex) begin
        counters_17 <= _T_7;
      end
    end
    if (reset) begin
      counters_18 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h12 == io_lastIndex) begin
            counters_18 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h12 == io_lastIndex) begin
            counters_18 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h12 == io_lastIndex) begin
          counters_18 <= _T_4;
        end
      end else if (5'h12 == io_lastIndex) begin
        counters_18 <= _T_7;
      end
    end
    if (reset) begin
      counters_19 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h13 == io_lastIndex) begin
            counters_19 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h13 == io_lastIndex) begin
            counters_19 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h13 == io_lastIndex) begin
          counters_19 <= _T_4;
        end
      end else if (5'h13 == io_lastIndex) begin
        counters_19 <= _T_7;
      end
    end
    if (reset) begin
      counters_20 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h14 == io_lastIndex) begin
            counters_20 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h14 == io_lastIndex) begin
            counters_20 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h14 == io_lastIndex) begin
          counters_20 <= _T_4;
        end
      end else if (5'h14 == io_lastIndex) begin
        counters_20 <= _T_7;
      end
    end
    if (reset) begin
      counters_21 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h15 == io_lastIndex) begin
            counters_21 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h15 == io_lastIndex) begin
            counters_21 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h15 == io_lastIndex) begin
          counters_21 <= _T_4;
        end
      end else if (5'h15 == io_lastIndex) begin
        counters_21 <= _T_7;
      end
    end
    if (reset) begin
      counters_22 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h16 == io_lastIndex) begin
            counters_22 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h16 == io_lastIndex) begin
            counters_22 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h16 == io_lastIndex) begin
          counters_22 <= _T_4;
        end
      end else if (5'h16 == io_lastIndex) begin
        counters_22 <= _T_7;
      end
    end
    if (reset) begin
      counters_23 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h17 == io_lastIndex) begin
            counters_23 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h17 == io_lastIndex) begin
            counters_23 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h17 == io_lastIndex) begin
          counters_23 <= _T_4;
        end
      end else if (5'h17 == io_lastIndex) begin
        counters_23 <= _T_7;
      end
    end
    if (reset) begin
      counters_24 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h18 == io_lastIndex) begin
            counters_24 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h18 == io_lastIndex) begin
            counters_24 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h18 == io_lastIndex) begin
          counters_24 <= _T_4;
        end
      end else if (5'h18 == io_lastIndex) begin
        counters_24 <= _T_7;
      end
    end
    if (reset) begin
      counters_25 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h19 == io_lastIndex) begin
            counters_25 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h19 == io_lastIndex) begin
            counters_25 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h19 == io_lastIndex) begin
          counters_25 <= _T_4;
        end
      end else if (5'h19 == io_lastIndex) begin
        counters_25 <= _T_7;
      end
    end
    if (reset) begin
      counters_26 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h1a == io_lastIndex) begin
            counters_26 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h1a == io_lastIndex) begin
            counters_26 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h1a == io_lastIndex) begin
          counters_26 <= _T_4;
        end
      end else if (5'h1a == io_lastIndex) begin
        counters_26 <= _T_7;
      end
    end
    if (reset) begin
      counters_27 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h1b == io_lastIndex) begin
            counters_27 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h1b == io_lastIndex) begin
            counters_27 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h1b == io_lastIndex) begin
          counters_27 <= _T_4;
        end
      end else if (5'h1b == io_lastIndex) begin
        counters_27 <= _T_7;
      end
    end
    if (reset) begin
      counters_28 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h1c == io_lastIndex) begin
            counters_28 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h1c == io_lastIndex) begin
            counters_28 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h1c == io_lastIndex) begin
          counters_28 <= _T_4;
        end
      end else if (5'h1c == io_lastIndex) begin
        counters_28 <= _T_7;
      end
    end
    if (reset) begin
      counters_29 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h1d == io_lastIndex) begin
            counters_29 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h1d == io_lastIndex) begin
            counters_29 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h1d == io_lastIndex) begin
          counters_29 <= _T_4;
        end
      end else if (5'h1d == io_lastIndex) begin
        counters_29 <= _T_7;
      end
    end
    if (reset) begin
      counters_30 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h1e == io_lastIndex) begin
            counters_30 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h1e == io_lastIndex) begin
            counters_30 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h1e == io_lastIndex) begin
          counters_30 <= _T_4;
        end
      end else if (5'h1e == io_lastIndex) begin
        counters_30 <= _T_7;
      end
    end
    if (reset) begin
      counters_31 <= 2'h2;
    end else if (io_lastBranch) begin
      if (_T_1) begin
        if (_T_2) begin
          if (5'h1f == io_lastIndex) begin
            counters_31 <= _T_4;
          end
        end
      end else if (_T_5) begin
        if (io_lastTaken) begin
          if (5'h1f == io_lastIndex) begin
            counters_31 <= _T_7;
          end
        end
      end else if (_T_2) begin
        if (5'h1f == io_lastIndex) begin
          counters_31 <= _T_4;
        end
      end else if (5'h1f == io_lastIndex) begin
        counters_31 <= _T_7;
      end
    end
  end
endmodule
module BTB(
  input         clock,
  input         reset,
  input         io_branch,
  input         io_jump,
  input  [31:0] io_pc,
  input  [31:0] io_target,
  input  [31:0] io_lookupPc,
  output        io_lookupBranch,
  output        io_lookupJump,
  output [31:0] io_lookupTarget
);
  reg  lines_jump [0:63]; // @[BTB.scala 33:20]
  reg [31:0] _RAND_0;
  wire  lines_jump__T_5_data; // @[BTB.scala 33:20]
  wire [5:0] lines_jump__T_5_addr; // @[BTB.scala 33:20]
  wire  lines_jump__T_7_data; // @[BTB.scala 33:20]
  wire [5:0] lines_jump__T_7_addr; // @[BTB.scala 33:20]
  wire  lines_jump__T_9_data; // @[BTB.scala 33:20]
  wire [5:0] lines_jump__T_9_addr; // @[BTB.scala 33:20]
  wire  lines_jump__T_1_data; // @[BTB.scala 33:20]
  wire [5:0] lines_jump__T_1_addr; // @[BTB.scala 33:20]
  wire  lines_jump__T_1_mask; // @[BTB.scala 33:20]
  wire  lines_jump__T_1_en; // @[BTB.scala 33:20]
  wire  lines_jump__T_2_data; // @[BTB.scala 33:20]
  wire [5:0] lines_jump__T_2_addr; // @[BTB.scala 33:20]
  wire  lines_jump__T_2_mask; // @[BTB.scala 33:20]
  wire  lines_jump__T_2_en; // @[BTB.scala 33:20]
  wire  lines_jump__T_3_data; // @[BTB.scala 33:20]
  wire [5:0] lines_jump__T_3_addr; // @[BTB.scala 33:20]
  wire  lines_jump__T_3_mask; // @[BTB.scala 33:20]
  wire  lines_jump__T_3_en; // @[BTB.scala 33:20]
  reg [23:0] lines_pc [0:63]; // @[BTB.scala 33:20]
  reg [31:0] _RAND_1;
  wire [23:0] lines_pc__T_5_data; // @[BTB.scala 33:20]
  wire [5:0] lines_pc__T_5_addr; // @[BTB.scala 33:20]
  wire [23:0] lines_pc__T_7_data; // @[BTB.scala 33:20]
  wire [5:0] lines_pc__T_7_addr; // @[BTB.scala 33:20]
  wire [23:0] lines_pc__T_9_data; // @[BTB.scala 33:20]
  wire [5:0] lines_pc__T_9_addr; // @[BTB.scala 33:20]
  wire [23:0] lines_pc__T_1_data; // @[BTB.scala 33:20]
  wire [5:0] lines_pc__T_1_addr; // @[BTB.scala 33:20]
  wire  lines_pc__T_1_mask; // @[BTB.scala 33:20]
  wire  lines_pc__T_1_en; // @[BTB.scala 33:20]
  wire [23:0] lines_pc__T_2_data; // @[BTB.scala 33:20]
  wire [5:0] lines_pc__T_2_addr; // @[BTB.scala 33:20]
  wire  lines_pc__T_2_mask; // @[BTB.scala 33:20]
  wire  lines_pc__T_2_en; // @[BTB.scala 33:20]
  wire [23:0] lines_pc__T_3_data; // @[BTB.scala 33:20]
  wire [5:0] lines_pc__T_3_addr; // @[BTB.scala 33:20]
  wire  lines_pc__T_3_mask; // @[BTB.scala 33:20]
  wire  lines_pc__T_3_en; // @[BTB.scala 33:20]
  reg [29:0] lines_target [0:63]; // @[BTB.scala 33:20]
  reg [31:0] _RAND_2;
  wire [29:0] lines_target__T_5_data; // @[BTB.scala 33:20]
  wire [5:0] lines_target__T_5_addr; // @[BTB.scala 33:20]
  wire [29:0] lines_target__T_7_data; // @[BTB.scala 33:20]
  wire [5:0] lines_target__T_7_addr; // @[BTB.scala 33:20]
  wire [29:0] lines_target__T_9_data; // @[BTB.scala 33:20]
  wire [5:0] lines_target__T_9_addr; // @[BTB.scala 33:20]
  wire [29:0] lines_target__T_1_data; // @[BTB.scala 33:20]
  wire [5:0] lines_target__T_1_addr; // @[BTB.scala 33:20]
  wire  lines_target__T_1_mask; // @[BTB.scala 33:20]
  wire  lines_target__T_1_en; // @[BTB.scala 33:20]
  wire [29:0] lines_target__T_2_data; // @[BTB.scala 33:20]
  wire [5:0] lines_target__T_2_addr; // @[BTB.scala 33:20]
  wire  lines_target__T_2_mask; // @[BTB.scala 33:20]
  wire  lines_target__T_2_en; // @[BTB.scala 33:20]
  wire [29:0] lines_target__T_3_data; // @[BTB.scala 33:20]
  wire [5:0] lines_target__T_3_addr; // @[BTB.scala 33:20]
  wire  lines_target__T_3_mask; // @[BTB.scala 33:20]
  wire  lines_target__T_3_en; // @[BTB.scala 33:20]
  reg  valids_0; // @[BTB.scala 32:24]
  reg [31:0] _RAND_3;
  reg  valids_1; // @[BTB.scala 32:24]
  reg [31:0] _RAND_4;
  reg  valids_2; // @[BTB.scala 32:24]
  reg [31:0] _RAND_5;
  reg  valids_3; // @[BTB.scala 32:24]
  reg [31:0] _RAND_6;
  reg  valids_4; // @[BTB.scala 32:24]
  reg [31:0] _RAND_7;
  reg  valids_5; // @[BTB.scala 32:24]
  reg [31:0] _RAND_8;
  reg  valids_6; // @[BTB.scala 32:24]
  reg [31:0] _RAND_9;
  reg  valids_7; // @[BTB.scala 32:24]
  reg [31:0] _RAND_10;
  reg  valids_8; // @[BTB.scala 32:24]
  reg [31:0] _RAND_11;
  reg  valids_9; // @[BTB.scala 32:24]
  reg [31:0] _RAND_12;
  reg  valids_10; // @[BTB.scala 32:24]
  reg [31:0] _RAND_13;
  reg  valids_11; // @[BTB.scala 32:24]
  reg [31:0] _RAND_14;
  reg  valids_12; // @[BTB.scala 32:24]
  reg [31:0] _RAND_15;
  reg  valids_13; // @[BTB.scala 32:24]
  reg [31:0] _RAND_16;
  reg  valids_14; // @[BTB.scala 32:24]
  reg [31:0] _RAND_17;
  reg  valids_15; // @[BTB.scala 32:24]
  reg [31:0] _RAND_18;
  reg  valids_16; // @[BTB.scala 32:24]
  reg [31:0] _RAND_19;
  reg  valids_17; // @[BTB.scala 32:24]
  reg [31:0] _RAND_20;
  reg  valids_18; // @[BTB.scala 32:24]
  reg [31:0] _RAND_21;
  reg  valids_19; // @[BTB.scala 32:24]
  reg [31:0] _RAND_22;
  reg  valids_20; // @[BTB.scala 32:24]
  reg [31:0] _RAND_23;
  reg  valids_21; // @[BTB.scala 32:24]
  reg [31:0] _RAND_24;
  reg  valids_22; // @[BTB.scala 32:24]
  reg [31:0] _RAND_25;
  reg  valids_23; // @[BTB.scala 32:24]
  reg [31:0] _RAND_26;
  reg  valids_24; // @[BTB.scala 32:24]
  reg [31:0] _RAND_27;
  reg  valids_25; // @[BTB.scala 32:24]
  reg [31:0] _RAND_28;
  reg  valids_26; // @[BTB.scala 32:24]
  reg [31:0] _RAND_29;
  reg  valids_27; // @[BTB.scala 32:24]
  reg [31:0] _RAND_30;
  reg  valids_28; // @[BTB.scala 32:24]
  reg [31:0] _RAND_31;
  reg  valids_29; // @[BTB.scala 32:24]
  reg [31:0] _RAND_32;
  reg  valids_30; // @[BTB.scala 32:24]
  reg [31:0] _RAND_33;
  reg  valids_31; // @[BTB.scala 32:24]
  reg [31:0] _RAND_34;
  reg  valids_32; // @[BTB.scala 32:24]
  reg [31:0] _RAND_35;
  reg  valids_33; // @[BTB.scala 32:24]
  reg [31:0] _RAND_36;
  reg  valids_34; // @[BTB.scala 32:24]
  reg [31:0] _RAND_37;
  reg  valids_35; // @[BTB.scala 32:24]
  reg [31:0] _RAND_38;
  reg  valids_36; // @[BTB.scala 32:24]
  reg [31:0] _RAND_39;
  reg  valids_37; // @[BTB.scala 32:24]
  reg [31:0] _RAND_40;
  reg  valids_38; // @[BTB.scala 32:24]
  reg [31:0] _RAND_41;
  reg  valids_39; // @[BTB.scala 32:24]
  reg [31:0] _RAND_42;
  reg  valids_40; // @[BTB.scala 32:24]
  reg [31:0] _RAND_43;
  reg  valids_41; // @[BTB.scala 32:24]
  reg [31:0] _RAND_44;
  reg  valids_42; // @[BTB.scala 32:24]
  reg [31:0] _RAND_45;
  reg  valids_43; // @[BTB.scala 32:24]
  reg [31:0] _RAND_46;
  reg  valids_44; // @[BTB.scala 32:24]
  reg [31:0] _RAND_47;
  reg  valids_45; // @[BTB.scala 32:24]
  reg [31:0] _RAND_48;
  reg  valids_46; // @[BTB.scala 32:24]
  reg [31:0] _RAND_49;
  reg  valids_47; // @[BTB.scala 32:24]
  reg [31:0] _RAND_50;
  reg  valids_48; // @[BTB.scala 32:24]
  reg [31:0] _RAND_51;
  reg  valids_49; // @[BTB.scala 32:24]
  reg [31:0] _RAND_52;
  reg  valids_50; // @[BTB.scala 32:24]
  reg [31:0] _RAND_53;
  reg  valids_51; // @[BTB.scala 32:24]
  reg [31:0] _RAND_54;
  reg  valids_52; // @[BTB.scala 32:24]
  reg [31:0] _RAND_55;
  reg  valids_53; // @[BTB.scala 32:24]
  reg [31:0] _RAND_56;
  reg  valids_54; // @[BTB.scala 32:24]
  reg [31:0] _RAND_57;
  reg  valids_55; // @[BTB.scala 32:24]
  reg [31:0] _RAND_58;
  reg  valids_56; // @[BTB.scala 32:24]
  reg [31:0] _RAND_59;
  reg  valids_57; // @[BTB.scala 32:24]
  reg [31:0] _RAND_60;
  reg  valids_58; // @[BTB.scala 32:24]
  reg [31:0] _RAND_61;
  reg  valids_59; // @[BTB.scala 32:24]
  reg [31:0] _RAND_62;
  reg  valids_60; // @[BTB.scala 32:24]
  reg [31:0] _RAND_63;
  reg  valids_61; // @[BTB.scala 32:24]
  reg [31:0] _RAND_64;
  reg  valids_62; // @[BTB.scala 32:24]
  reg [31:0] _RAND_65;
  reg  valids_63; // @[BTB.scala 32:24]
  reg [31:0] _RAND_66;
  wire [5:0] index = io_pc[7:2]; // @[BTB.scala 36:22]
  wire  _GEN_200 = 6'h0 == index; // @[BTB.scala 42:25]
  wire  _GEN_0 = _GEN_200 | valids_0; // @[BTB.scala 42:25]
  wire  _GEN_201 = 6'h1 == index; // @[BTB.scala 42:25]
  wire  _GEN_1 = _GEN_201 | valids_1; // @[BTB.scala 42:25]
  wire  _GEN_202 = 6'h2 == index; // @[BTB.scala 42:25]
  wire  _GEN_2 = _GEN_202 | valids_2; // @[BTB.scala 42:25]
  wire  _GEN_203 = 6'h3 == index; // @[BTB.scala 42:25]
  wire  _GEN_3 = _GEN_203 | valids_3; // @[BTB.scala 42:25]
  wire  _GEN_204 = 6'h4 == index; // @[BTB.scala 42:25]
  wire  _GEN_4 = _GEN_204 | valids_4; // @[BTB.scala 42:25]
  wire  _GEN_205 = 6'h5 == index; // @[BTB.scala 42:25]
  wire  _GEN_5 = _GEN_205 | valids_5; // @[BTB.scala 42:25]
  wire  _GEN_206 = 6'h6 == index; // @[BTB.scala 42:25]
  wire  _GEN_6 = _GEN_206 | valids_6; // @[BTB.scala 42:25]
  wire  _GEN_207 = 6'h7 == index; // @[BTB.scala 42:25]
  wire  _GEN_7 = _GEN_207 | valids_7; // @[BTB.scala 42:25]
  wire  _GEN_208 = 6'h8 == index; // @[BTB.scala 42:25]
  wire  _GEN_8 = _GEN_208 | valids_8; // @[BTB.scala 42:25]
  wire  _GEN_209 = 6'h9 == index; // @[BTB.scala 42:25]
  wire  _GEN_9 = _GEN_209 | valids_9; // @[BTB.scala 42:25]
  wire  _GEN_210 = 6'ha == index; // @[BTB.scala 42:25]
  wire  _GEN_10 = _GEN_210 | valids_10; // @[BTB.scala 42:25]
  wire  _GEN_211 = 6'hb == index; // @[BTB.scala 42:25]
  wire  _GEN_11 = _GEN_211 | valids_11; // @[BTB.scala 42:25]
  wire  _GEN_212 = 6'hc == index; // @[BTB.scala 42:25]
  wire  _GEN_12 = _GEN_212 | valids_12; // @[BTB.scala 42:25]
  wire  _GEN_213 = 6'hd == index; // @[BTB.scala 42:25]
  wire  _GEN_13 = _GEN_213 | valids_13; // @[BTB.scala 42:25]
  wire  _GEN_214 = 6'he == index; // @[BTB.scala 42:25]
  wire  _GEN_14 = _GEN_214 | valids_14; // @[BTB.scala 42:25]
  wire  _GEN_215 = 6'hf == index; // @[BTB.scala 42:25]
  wire  _GEN_15 = _GEN_215 | valids_15; // @[BTB.scala 42:25]
  wire  _GEN_216 = 6'h10 == index; // @[BTB.scala 42:25]
  wire  _GEN_16 = _GEN_216 | valids_16; // @[BTB.scala 42:25]
  wire  _GEN_217 = 6'h11 == index; // @[BTB.scala 42:25]
  wire  _GEN_17 = _GEN_217 | valids_17; // @[BTB.scala 42:25]
  wire  _GEN_218 = 6'h12 == index; // @[BTB.scala 42:25]
  wire  _GEN_18 = _GEN_218 | valids_18; // @[BTB.scala 42:25]
  wire  _GEN_219 = 6'h13 == index; // @[BTB.scala 42:25]
  wire  _GEN_19 = _GEN_219 | valids_19; // @[BTB.scala 42:25]
  wire  _GEN_220 = 6'h14 == index; // @[BTB.scala 42:25]
  wire  _GEN_20 = _GEN_220 | valids_20; // @[BTB.scala 42:25]
  wire  _GEN_221 = 6'h15 == index; // @[BTB.scala 42:25]
  wire  _GEN_21 = _GEN_221 | valids_21; // @[BTB.scala 42:25]
  wire  _GEN_222 = 6'h16 == index; // @[BTB.scala 42:25]
  wire  _GEN_22 = _GEN_222 | valids_22; // @[BTB.scala 42:25]
  wire  _GEN_223 = 6'h17 == index; // @[BTB.scala 42:25]
  wire  _GEN_23 = _GEN_223 | valids_23; // @[BTB.scala 42:25]
  wire  _GEN_224 = 6'h18 == index; // @[BTB.scala 42:25]
  wire  _GEN_24 = _GEN_224 | valids_24; // @[BTB.scala 42:25]
  wire  _GEN_225 = 6'h19 == index; // @[BTB.scala 42:25]
  wire  _GEN_25 = _GEN_225 | valids_25; // @[BTB.scala 42:25]
  wire  _GEN_226 = 6'h1a == index; // @[BTB.scala 42:25]
  wire  _GEN_26 = _GEN_226 | valids_26; // @[BTB.scala 42:25]
  wire  _GEN_227 = 6'h1b == index; // @[BTB.scala 42:25]
  wire  _GEN_27 = _GEN_227 | valids_27; // @[BTB.scala 42:25]
  wire  _GEN_228 = 6'h1c == index; // @[BTB.scala 42:25]
  wire  _GEN_28 = _GEN_228 | valids_28; // @[BTB.scala 42:25]
  wire  _GEN_229 = 6'h1d == index; // @[BTB.scala 42:25]
  wire  _GEN_29 = _GEN_229 | valids_29; // @[BTB.scala 42:25]
  wire  _GEN_230 = 6'h1e == index; // @[BTB.scala 42:25]
  wire  _GEN_30 = _GEN_230 | valids_30; // @[BTB.scala 42:25]
  wire  _GEN_231 = 6'h1f == index; // @[BTB.scala 42:25]
  wire  _GEN_31 = _GEN_231 | valids_31; // @[BTB.scala 42:25]
  wire  _GEN_232 = 6'h20 == index; // @[BTB.scala 42:25]
  wire  _GEN_32 = _GEN_232 | valids_32; // @[BTB.scala 42:25]
  wire  _GEN_233 = 6'h21 == index; // @[BTB.scala 42:25]
  wire  _GEN_33 = _GEN_233 | valids_33; // @[BTB.scala 42:25]
  wire  _GEN_234 = 6'h22 == index; // @[BTB.scala 42:25]
  wire  _GEN_34 = _GEN_234 | valids_34; // @[BTB.scala 42:25]
  wire  _GEN_235 = 6'h23 == index; // @[BTB.scala 42:25]
  wire  _GEN_35 = _GEN_235 | valids_35; // @[BTB.scala 42:25]
  wire  _GEN_236 = 6'h24 == index; // @[BTB.scala 42:25]
  wire  _GEN_36 = _GEN_236 | valids_36; // @[BTB.scala 42:25]
  wire  _GEN_237 = 6'h25 == index; // @[BTB.scala 42:25]
  wire  _GEN_37 = _GEN_237 | valids_37; // @[BTB.scala 42:25]
  wire  _GEN_238 = 6'h26 == index; // @[BTB.scala 42:25]
  wire  _GEN_38 = _GEN_238 | valids_38; // @[BTB.scala 42:25]
  wire  _GEN_239 = 6'h27 == index; // @[BTB.scala 42:25]
  wire  _GEN_39 = _GEN_239 | valids_39; // @[BTB.scala 42:25]
  wire  _GEN_240 = 6'h28 == index; // @[BTB.scala 42:25]
  wire  _GEN_40 = _GEN_240 | valids_40; // @[BTB.scala 42:25]
  wire  _GEN_241 = 6'h29 == index; // @[BTB.scala 42:25]
  wire  _GEN_41 = _GEN_241 | valids_41; // @[BTB.scala 42:25]
  wire  _GEN_242 = 6'h2a == index; // @[BTB.scala 42:25]
  wire  _GEN_42 = _GEN_242 | valids_42; // @[BTB.scala 42:25]
  wire  _GEN_243 = 6'h2b == index; // @[BTB.scala 42:25]
  wire  _GEN_43 = _GEN_243 | valids_43; // @[BTB.scala 42:25]
  wire  _GEN_244 = 6'h2c == index; // @[BTB.scala 42:25]
  wire  _GEN_44 = _GEN_244 | valids_44; // @[BTB.scala 42:25]
  wire  _GEN_245 = 6'h2d == index; // @[BTB.scala 42:25]
  wire  _GEN_45 = _GEN_245 | valids_45; // @[BTB.scala 42:25]
  wire  _GEN_246 = 6'h2e == index; // @[BTB.scala 42:25]
  wire  _GEN_46 = _GEN_246 | valids_46; // @[BTB.scala 42:25]
  wire  _GEN_247 = 6'h2f == index; // @[BTB.scala 42:25]
  wire  _GEN_47 = _GEN_247 | valids_47; // @[BTB.scala 42:25]
  wire  _GEN_248 = 6'h30 == index; // @[BTB.scala 42:25]
  wire  _GEN_48 = _GEN_248 | valids_48; // @[BTB.scala 42:25]
  wire  _GEN_249 = 6'h31 == index; // @[BTB.scala 42:25]
  wire  _GEN_49 = _GEN_249 | valids_49; // @[BTB.scala 42:25]
  wire  _GEN_250 = 6'h32 == index; // @[BTB.scala 42:25]
  wire  _GEN_50 = _GEN_250 | valids_50; // @[BTB.scala 42:25]
  wire  _GEN_251 = 6'h33 == index; // @[BTB.scala 42:25]
  wire  _GEN_51 = _GEN_251 | valids_51; // @[BTB.scala 42:25]
  wire  _GEN_252 = 6'h34 == index; // @[BTB.scala 42:25]
  wire  _GEN_52 = _GEN_252 | valids_52; // @[BTB.scala 42:25]
  wire  _GEN_253 = 6'h35 == index; // @[BTB.scala 42:25]
  wire  _GEN_53 = _GEN_253 | valids_53; // @[BTB.scala 42:25]
  wire  _GEN_254 = 6'h36 == index; // @[BTB.scala 42:25]
  wire  _GEN_54 = _GEN_254 | valids_54; // @[BTB.scala 42:25]
  wire  _GEN_255 = 6'h37 == index; // @[BTB.scala 42:25]
  wire  _GEN_55 = _GEN_255 | valids_55; // @[BTB.scala 42:25]
  wire  _GEN_256 = 6'h38 == index; // @[BTB.scala 42:25]
  wire  _GEN_56 = _GEN_256 | valids_56; // @[BTB.scala 42:25]
  wire  _GEN_257 = 6'h39 == index; // @[BTB.scala 42:25]
  wire  _GEN_57 = _GEN_257 | valids_57; // @[BTB.scala 42:25]
  wire  _GEN_258 = 6'h3a == index; // @[BTB.scala 42:25]
  wire  _GEN_58 = _GEN_258 | valids_58; // @[BTB.scala 42:25]
  wire  _GEN_259 = 6'h3b == index; // @[BTB.scala 42:25]
  wire  _GEN_59 = _GEN_259 | valids_59; // @[BTB.scala 42:25]
  wire  _GEN_260 = 6'h3c == index; // @[BTB.scala 42:25]
  wire  _GEN_60 = _GEN_260 | valids_60; // @[BTB.scala 42:25]
  wire  _GEN_261 = 6'h3d == index; // @[BTB.scala 42:25]
  wire  _GEN_61 = _GEN_261 | valids_61; // @[BTB.scala 42:25]
  wire  _GEN_262 = 6'h3e == index; // @[BTB.scala 42:25]
  wire  _GEN_62 = _GEN_262 | valids_62; // @[BTB.scala 42:25]
  wire  _GEN_263 = 6'h3f == index; // @[BTB.scala 42:25]
  wire  _GEN_63 = _GEN_263 | valids_63; // @[BTB.scala 42:25]
  wire [5:0] lookupIndex = io_lookupPc[7:2]; // @[BTB.scala 49:32]
  wire [23:0] lookupPcSel = io_lookupPc[31:8]; // @[BTB.scala 51:32]
  wire  _T_6 = lines_pc__T_5_data == lookupPcSel; // @[BTB.scala 54:43]
  wire  _GEN_137 = 6'h1 == lookupIndex ? valids_1 : valids_0; // @[BTB.scala 53:41]
  wire  _GEN_138 = 6'h2 == lookupIndex ? valids_2 : _GEN_137; // @[BTB.scala 53:41]
  wire  _GEN_139 = 6'h3 == lookupIndex ? valids_3 : _GEN_138; // @[BTB.scala 53:41]
  wire  _GEN_140 = 6'h4 == lookupIndex ? valids_4 : _GEN_139; // @[BTB.scala 53:41]
  wire  _GEN_141 = 6'h5 == lookupIndex ? valids_5 : _GEN_140; // @[BTB.scala 53:41]
  wire  _GEN_142 = 6'h6 == lookupIndex ? valids_6 : _GEN_141; // @[BTB.scala 53:41]
  wire  _GEN_143 = 6'h7 == lookupIndex ? valids_7 : _GEN_142; // @[BTB.scala 53:41]
  wire  _GEN_144 = 6'h8 == lookupIndex ? valids_8 : _GEN_143; // @[BTB.scala 53:41]
  wire  _GEN_145 = 6'h9 == lookupIndex ? valids_9 : _GEN_144; // @[BTB.scala 53:41]
  wire  _GEN_146 = 6'ha == lookupIndex ? valids_10 : _GEN_145; // @[BTB.scala 53:41]
  wire  _GEN_147 = 6'hb == lookupIndex ? valids_11 : _GEN_146; // @[BTB.scala 53:41]
  wire  _GEN_148 = 6'hc == lookupIndex ? valids_12 : _GEN_147; // @[BTB.scala 53:41]
  wire  _GEN_149 = 6'hd == lookupIndex ? valids_13 : _GEN_148; // @[BTB.scala 53:41]
  wire  _GEN_150 = 6'he == lookupIndex ? valids_14 : _GEN_149; // @[BTB.scala 53:41]
  wire  _GEN_151 = 6'hf == lookupIndex ? valids_15 : _GEN_150; // @[BTB.scala 53:41]
  wire  _GEN_152 = 6'h10 == lookupIndex ? valids_16 : _GEN_151; // @[BTB.scala 53:41]
  wire  _GEN_153 = 6'h11 == lookupIndex ? valids_17 : _GEN_152; // @[BTB.scala 53:41]
  wire  _GEN_154 = 6'h12 == lookupIndex ? valids_18 : _GEN_153; // @[BTB.scala 53:41]
  wire  _GEN_155 = 6'h13 == lookupIndex ? valids_19 : _GEN_154; // @[BTB.scala 53:41]
  wire  _GEN_156 = 6'h14 == lookupIndex ? valids_20 : _GEN_155; // @[BTB.scala 53:41]
  wire  _GEN_157 = 6'h15 == lookupIndex ? valids_21 : _GEN_156; // @[BTB.scala 53:41]
  wire  _GEN_158 = 6'h16 == lookupIndex ? valids_22 : _GEN_157; // @[BTB.scala 53:41]
  wire  _GEN_159 = 6'h17 == lookupIndex ? valids_23 : _GEN_158; // @[BTB.scala 53:41]
  wire  _GEN_160 = 6'h18 == lookupIndex ? valids_24 : _GEN_159; // @[BTB.scala 53:41]
  wire  _GEN_161 = 6'h19 == lookupIndex ? valids_25 : _GEN_160; // @[BTB.scala 53:41]
  wire  _GEN_162 = 6'h1a == lookupIndex ? valids_26 : _GEN_161; // @[BTB.scala 53:41]
  wire  _GEN_163 = 6'h1b == lookupIndex ? valids_27 : _GEN_162; // @[BTB.scala 53:41]
  wire  _GEN_164 = 6'h1c == lookupIndex ? valids_28 : _GEN_163; // @[BTB.scala 53:41]
  wire  _GEN_165 = 6'h1d == lookupIndex ? valids_29 : _GEN_164; // @[BTB.scala 53:41]
  wire  _GEN_166 = 6'h1e == lookupIndex ? valids_30 : _GEN_165; // @[BTB.scala 53:41]
  wire  _GEN_167 = 6'h1f == lookupIndex ? valids_31 : _GEN_166; // @[BTB.scala 53:41]
  wire  _GEN_168 = 6'h20 == lookupIndex ? valids_32 : _GEN_167; // @[BTB.scala 53:41]
  wire  _GEN_169 = 6'h21 == lookupIndex ? valids_33 : _GEN_168; // @[BTB.scala 53:41]
  wire  _GEN_170 = 6'h22 == lookupIndex ? valids_34 : _GEN_169; // @[BTB.scala 53:41]
  wire  _GEN_171 = 6'h23 == lookupIndex ? valids_35 : _GEN_170; // @[BTB.scala 53:41]
  wire  _GEN_172 = 6'h24 == lookupIndex ? valids_36 : _GEN_171; // @[BTB.scala 53:41]
  wire  _GEN_173 = 6'h25 == lookupIndex ? valids_37 : _GEN_172; // @[BTB.scala 53:41]
  wire  _GEN_174 = 6'h26 == lookupIndex ? valids_38 : _GEN_173; // @[BTB.scala 53:41]
  wire  _GEN_175 = 6'h27 == lookupIndex ? valids_39 : _GEN_174; // @[BTB.scala 53:41]
  wire  _GEN_176 = 6'h28 == lookupIndex ? valids_40 : _GEN_175; // @[BTB.scala 53:41]
  wire  _GEN_177 = 6'h29 == lookupIndex ? valids_41 : _GEN_176; // @[BTB.scala 53:41]
  wire  _GEN_178 = 6'h2a == lookupIndex ? valids_42 : _GEN_177; // @[BTB.scala 53:41]
  wire  _GEN_179 = 6'h2b == lookupIndex ? valids_43 : _GEN_178; // @[BTB.scala 53:41]
  wire  _GEN_180 = 6'h2c == lookupIndex ? valids_44 : _GEN_179; // @[BTB.scala 53:41]
  wire  _GEN_181 = 6'h2d == lookupIndex ? valids_45 : _GEN_180; // @[BTB.scala 53:41]
  wire  _GEN_182 = 6'h2e == lookupIndex ? valids_46 : _GEN_181; // @[BTB.scala 53:41]
  wire  _GEN_183 = 6'h2f == lookupIndex ? valids_47 : _GEN_182; // @[BTB.scala 53:41]
  wire  _GEN_184 = 6'h30 == lookupIndex ? valids_48 : _GEN_183; // @[BTB.scala 53:41]
  wire  _GEN_185 = 6'h31 == lookupIndex ? valids_49 : _GEN_184; // @[BTB.scala 53:41]
  wire  _GEN_186 = 6'h32 == lookupIndex ? valids_50 : _GEN_185; // @[BTB.scala 53:41]
  wire  _GEN_187 = 6'h33 == lookupIndex ? valids_51 : _GEN_186; // @[BTB.scala 53:41]
  wire  _GEN_188 = 6'h34 == lookupIndex ? valids_52 : _GEN_187; // @[BTB.scala 53:41]
  wire  _GEN_189 = 6'h35 == lookupIndex ? valids_53 : _GEN_188; // @[BTB.scala 53:41]
  wire  _GEN_190 = 6'h36 == lookupIndex ? valids_54 : _GEN_189; // @[BTB.scala 53:41]
  wire  _GEN_191 = 6'h37 == lookupIndex ? valids_55 : _GEN_190; // @[BTB.scala 53:41]
  wire  _GEN_192 = 6'h38 == lookupIndex ? valids_56 : _GEN_191; // @[BTB.scala 53:41]
  wire  _GEN_193 = 6'h39 == lookupIndex ? valids_57 : _GEN_192; // @[BTB.scala 53:41]
  wire  _GEN_194 = 6'h3a == lookupIndex ? valids_58 : _GEN_193; // @[BTB.scala 53:41]
  wire  _GEN_195 = 6'h3b == lookupIndex ? valids_59 : _GEN_194; // @[BTB.scala 53:41]
  wire  _GEN_196 = 6'h3c == lookupIndex ? valids_60 : _GEN_195; // @[BTB.scala 53:41]
  wire  _GEN_197 = 6'h3d == lookupIndex ? valids_61 : _GEN_196; // @[BTB.scala 53:41]
  wire  _GEN_198 = 6'h3e == lookupIndex ? valids_62 : _GEN_197; // @[BTB.scala 53:41]
  wire  _GEN_199 = 6'h3f == lookupIndex ? valids_63 : _GEN_198; // @[BTB.scala 53:41]
  wire  btbHit = _GEN_199 & _T_6; // @[BTB.scala 53:41]
  wire [29:0] _T_10 = btbHit ? lines_target__T_9_data : 30'h0; // @[BTB.scala 59:29]
  assign lines_jump__T_5_addr = io_lookupPc[7:2];
  assign lines_jump__T_5_data = lines_jump[lines_jump__T_5_addr]; // @[BTB.scala 33:20]
  assign lines_jump__T_7_addr = io_lookupPc[7:2];
  assign lines_jump__T_7_data = lines_jump[lines_jump__T_7_addr]; // @[BTB.scala 33:20]
  assign lines_jump__T_9_addr = io_lookupPc[7:2];
  assign lines_jump__T_9_data = lines_jump[lines_jump__T_9_addr]; // @[BTB.scala 33:20]
  assign lines_jump__T_1_data = io_jump;
  assign lines_jump__T_1_addr = io_pc[7:2];
  assign lines_jump__T_1_mask = 1'h1;
  assign lines_jump__T_1_en = io_branch;
  assign lines_jump__T_2_data = 1'h0;
  assign lines_jump__T_2_addr = io_pc[7:2];
  assign lines_jump__T_2_mask = 1'h0;
  assign lines_jump__T_2_en = io_branch;
  assign lines_jump__T_3_data = 1'h0;
  assign lines_jump__T_3_addr = io_pc[7:2];
  assign lines_jump__T_3_mask = 1'h0;
  assign lines_jump__T_3_en = io_branch;
  assign lines_pc__T_5_addr = io_lookupPc[7:2];
  assign lines_pc__T_5_data = lines_pc[lines_pc__T_5_addr]; // @[BTB.scala 33:20]
  assign lines_pc__T_7_addr = io_lookupPc[7:2];
  assign lines_pc__T_7_data = lines_pc[lines_pc__T_7_addr]; // @[BTB.scala 33:20]
  assign lines_pc__T_9_addr = io_lookupPc[7:2];
  assign lines_pc__T_9_data = lines_pc[lines_pc__T_9_addr]; // @[BTB.scala 33:20]
  assign lines_pc__T_1_data = 24'h0;
  assign lines_pc__T_1_addr = io_pc[7:2];
  assign lines_pc__T_1_mask = 1'h0;
  assign lines_pc__T_1_en = io_branch;
  assign lines_pc__T_2_data = io_pc[31:8];
  assign lines_pc__T_2_addr = io_pc[7:2];
  assign lines_pc__T_2_mask = 1'h1;
  assign lines_pc__T_2_en = io_branch;
  assign lines_pc__T_3_data = 24'h0;
  assign lines_pc__T_3_addr = io_pc[7:2];
  assign lines_pc__T_3_mask = 1'h0;
  assign lines_pc__T_3_en = io_branch;
  assign lines_target__T_5_addr = io_lookupPc[7:2];
  assign lines_target__T_5_data = lines_target[lines_target__T_5_addr]; // @[BTB.scala 33:20]
  assign lines_target__T_7_addr = io_lookupPc[7:2];
  assign lines_target__T_7_data = lines_target[lines_target__T_7_addr]; // @[BTB.scala 33:20]
  assign lines_target__T_9_addr = io_lookupPc[7:2];
  assign lines_target__T_9_data = lines_target[lines_target__T_9_addr]; // @[BTB.scala 33:20]
  assign lines_target__T_1_data = 30'h0;
  assign lines_target__T_1_addr = io_pc[7:2];
  assign lines_target__T_1_mask = 1'h0;
  assign lines_target__T_1_en = io_branch;
  assign lines_target__T_2_data = 30'h0;
  assign lines_target__T_2_addr = io_pc[7:2];
  assign lines_target__T_2_mask = 1'h0;
  assign lines_target__T_2_en = io_branch;
  assign lines_target__T_3_data = io_target[31:2];
  assign lines_target__T_3_addr = io_pc[7:2];
  assign lines_target__T_3_mask = 1'h1;
  assign lines_target__T_3_en = io_branch;
  assign io_lookupBranch = _GEN_199 & _T_6; // @[BTB.scala 57:19]
  assign io_lookupJump = btbHit & lines_jump__T_7_data; // @[BTB.scala 58:19]
  assign io_lookupTarget = {_T_10,2'h0}; // @[BTB.scala 59:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    lines_jump[initvar] = _RAND_0[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    lines_pc[initvar] = _RAND_1[23:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    lines_target[initvar] = _RAND_2[29:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  valids_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  valids_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  valids_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  valids_3 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  valids_4 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  valids_5 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  valids_6 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  valids_7 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  valids_8 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  valids_9 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  valids_10 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  valids_11 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  valids_12 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  valids_13 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  valids_14 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  valids_15 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  valids_16 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valids_17 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  valids_18 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  valids_19 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  valids_20 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  valids_21 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  valids_22 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  valids_23 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  valids_24 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  valids_25 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  valids_26 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  valids_27 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  valids_28 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  valids_29 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  valids_30 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  valids_31 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  valids_32 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  valids_33 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  valids_34 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  valids_35 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  valids_36 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  valids_37 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  valids_38 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  valids_39 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  valids_40 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  valids_41 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  valids_42 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  valids_43 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  valids_44 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  valids_45 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  valids_46 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  valids_47 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  valids_48 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  valids_49 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  valids_50 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  valids_51 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  valids_52 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  valids_53 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  valids_54 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  valids_55 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  valids_56 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  valids_57 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  valids_58 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  valids_59 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  valids_60 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  valids_61 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  valids_62 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  valids_63 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(lines_jump__T_1_en & lines_jump__T_1_mask) begin
      lines_jump[lines_jump__T_1_addr] <= lines_jump__T_1_data; // @[BTB.scala 33:20]
    end
    if(lines_jump__T_2_en & lines_jump__T_2_mask) begin
      lines_jump[lines_jump__T_2_addr] <= lines_jump__T_2_data; // @[BTB.scala 33:20]
    end
    if(lines_jump__T_3_en & lines_jump__T_3_mask) begin
      lines_jump[lines_jump__T_3_addr] <= lines_jump__T_3_data; // @[BTB.scala 33:20]
    end
    if(lines_pc__T_1_en & lines_pc__T_1_mask) begin
      lines_pc[lines_pc__T_1_addr] <= lines_pc__T_1_data; // @[BTB.scala 33:20]
    end
    if(lines_pc__T_2_en & lines_pc__T_2_mask) begin
      lines_pc[lines_pc__T_2_addr] <= lines_pc__T_2_data; // @[BTB.scala 33:20]
    end
    if(lines_pc__T_3_en & lines_pc__T_3_mask) begin
      lines_pc[lines_pc__T_3_addr] <= lines_pc__T_3_data; // @[BTB.scala 33:20]
    end
    if(lines_target__T_1_en & lines_target__T_1_mask) begin
      lines_target[lines_target__T_1_addr] <= lines_target__T_1_data; // @[BTB.scala 33:20]
    end
    if(lines_target__T_2_en & lines_target__T_2_mask) begin
      lines_target[lines_target__T_2_addr] <= lines_target__T_2_data; // @[BTB.scala 33:20]
    end
    if(lines_target__T_3_en & lines_target__T_3_mask) begin
      lines_target[lines_target__T_3_addr] <= lines_target__T_3_data; // @[BTB.scala 33:20]
    end
    if (reset) begin
      valids_0 <= 1'h0;
    end else if (io_branch) begin
      valids_0 <= _GEN_0;
    end
    if (reset) begin
      valids_1 <= 1'h0;
    end else if (io_branch) begin
      valids_1 <= _GEN_1;
    end
    if (reset) begin
      valids_2 <= 1'h0;
    end else if (io_branch) begin
      valids_2 <= _GEN_2;
    end
    if (reset) begin
      valids_3 <= 1'h0;
    end else if (io_branch) begin
      valids_3 <= _GEN_3;
    end
    if (reset) begin
      valids_4 <= 1'h0;
    end else if (io_branch) begin
      valids_4 <= _GEN_4;
    end
    if (reset) begin
      valids_5 <= 1'h0;
    end else if (io_branch) begin
      valids_5 <= _GEN_5;
    end
    if (reset) begin
      valids_6 <= 1'h0;
    end else if (io_branch) begin
      valids_6 <= _GEN_6;
    end
    if (reset) begin
      valids_7 <= 1'h0;
    end else if (io_branch) begin
      valids_7 <= _GEN_7;
    end
    if (reset) begin
      valids_8 <= 1'h0;
    end else if (io_branch) begin
      valids_8 <= _GEN_8;
    end
    if (reset) begin
      valids_9 <= 1'h0;
    end else if (io_branch) begin
      valids_9 <= _GEN_9;
    end
    if (reset) begin
      valids_10 <= 1'h0;
    end else if (io_branch) begin
      valids_10 <= _GEN_10;
    end
    if (reset) begin
      valids_11 <= 1'h0;
    end else if (io_branch) begin
      valids_11 <= _GEN_11;
    end
    if (reset) begin
      valids_12 <= 1'h0;
    end else if (io_branch) begin
      valids_12 <= _GEN_12;
    end
    if (reset) begin
      valids_13 <= 1'h0;
    end else if (io_branch) begin
      valids_13 <= _GEN_13;
    end
    if (reset) begin
      valids_14 <= 1'h0;
    end else if (io_branch) begin
      valids_14 <= _GEN_14;
    end
    if (reset) begin
      valids_15 <= 1'h0;
    end else if (io_branch) begin
      valids_15 <= _GEN_15;
    end
    if (reset) begin
      valids_16 <= 1'h0;
    end else if (io_branch) begin
      valids_16 <= _GEN_16;
    end
    if (reset) begin
      valids_17 <= 1'h0;
    end else if (io_branch) begin
      valids_17 <= _GEN_17;
    end
    if (reset) begin
      valids_18 <= 1'h0;
    end else if (io_branch) begin
      valids_18 <= _GEN_18;
    end
    if (reset) begin
      valids_19 <= 1'h0;
    end else if (io_branch) begin
      valids_19 <= _GEN_19;
    end
    if (reset) begin
      valids_20 <= 1'h0;
    end else if (io_branch) begin
      valids_20 <= _GEN_20;
    end
    if (reset) begin
      valids_21 <= 1'h0;
    end else if (io_branch) begin
      valids_21 <= _GEN_21;
    end
    if (reset) begin
      valids_22 <= 1'h0;
    end else if (io_branch) begin
      valids_22 <= _GEN_22;
    end
    if (reset) begin
      valids_23 <= 1'h0;
    end else if (io_branch) begin
      valids_23 <= _GEN_23;
    end
    if (reset) begin
      valids_24 <= 1'h0;
    end else if (io_branch) begin
      valids_24 <= _GEN_24;
    end
    if (reset) begin
      valids_25 <= 1'h0;
    end else if (io_branch) begin
      valids_25 <= _GEN_25;
    end
    if (reset) begin
      valids_26 <= 1'h0;
    end else if (io_branch) begin
      valids_26 <= _GEN_26;
    end
    if (reset) begin
      valids_27 <= 1'h0;
    end else if (io_branch) begin
      valids_27 <= _GEN_27;
    end
    if (reset) begin
      valids_28 <= 1'h0;
    end else if (io_branch) begin
      valids_28 <= _GEN_28;
    end
    if (reset) begin
      valids_29 <= 1'h0;
    end else if (io_branch) begin
      valids_29 <= _GEN_29;
    end
    if (reset) begin
      valids_30 <= 1'h0;
    end else if (io_branch) begin
      valids_30 <= _GEN_30;
    end
    if (reset) begin
      valids_31 <= 1'h0;
    end else if (io_branch) begin
      valids_31 <= _GEN_31;
    end
    if (reset) begin
      valids_32 <= 1'h0;
    end else if (io_branch) begin
      valids_32 <= _GEN_32;
    end
    if (reset) begin
      valids_33 <= 1'h0;
    end else if (io_branch) begin
      valids_33 <= _GEN_33;
    end
    if (reset) begin
      valids_34 <= 1'h0;
    end else if (io_branch) begin
      valids_34 <= _GEN_34;
    end
    if (reset) begin
      valids_35 <= 1'h0;
    end else if (io_branch) begin
      valids_35 <= _GEN_35;
    end
    if (reset) begin
      valids_36 <= 1'h0;
    end else if (io_branch) begin
      valids_36 <= _GEN_36;
    end
    if (reset) begin
      valids_37 <= 1'h0;
    end else if (io_branch) begin
      valids_37 <= _GEN_37;
    end
    if (reset) begin
      valids_38 <= 1'h0;
    end else if (io_branch) begin
      valids_38 <= _GEN_38;
    end
    if (reset) begin
      valids_39 <= 1'h0;
    end else if (io_branch) begin
      valids_39 <= _GEN_39;
    end
    if (reset) begin
      valids_40 <= 1'h0;
    end else if (io_branch) begin
      valids_40 <= _GEN_40;
    end
    if (reset) begin
      valids_41 <= 1'h0;
    end else if (io_branch) begin
      valids_41 <= _GEN_41;
    end
    if (reset) begin
      valids_42 <= 1'h0;
    end else if (io_branch) begin
      valids_42 <= _GEN_42;
    end
    if (reset) begin
      valids_43 <= 1'h0;
    end else if (io_branch) begin
      valids_43 <= _GEN_43;
    end
    if (reset) begin
      valids_44 <= 1'h0;
    end else if (io_branch) begin
      valids_44 <= _GEN_44;
    end
    if (reset) begin
      valids_45 <= 1'h0;
    end else if (io_branch) begin
      valids_45 <= _GEN_45;
    end
    if (reset) begin
      valids_46 <= 1'h0;
    end else if (io_branch) begin
      valids_46 <= _GEN_46;
    end
    if (reset) begin
      valids_47 <= 1'h0;
    end else if (io_branch) begin
      valids_47 <= _GEN_47;
    end
    if (reset) begin
      valids_48 <= 1'h0;
    end else if (io_branch) begin
      valids_48 <= _GEN_48;
    end
    if (reset) begin
      valids_49 <= 1'h0;
    end else if (io_branch) begin
      valids_49 <= _GEN_49;
    end
    if (reset) begin
      valids_50 <= 1'h0;
    end else if (io_branch) begin
      valids_50 <= _GEN_50;
    end
    if (reset) begin
      valids_51 <= 1'h0;
    end else if (io_branch) begin
      valids_51 <= _GEN_51;
    end
    if (reset) begin
      valids_52 <= 1'h0;
    end else if (io_branch) begin
      valids_52 <= _GEN_52;
    end
    if (reset) begin
      valids_53 <= 1'h0;
    end else if (io_branch) begin
      valids_53 <= _GEN_53;
    end
    if (reset) begin
      valids_54 <= 1'h0;
    end else if (io_branch) begin
      valids_54 <= _GEN_54;
    end
    if (reset) begin
      valids_55 <= 1'h0;
    end else if (io_branch) begin
      valids_55 <= _GEN_55;
    end
    if (reset) begin
      valids_56 <= 1'h0;
    end else if (io_branch) begin
      valids_56 <= _GEN_56;
    end
    if (reset) begin
      valids_57 <= 1'h0;
    end else if (io_branch) begin
      valids_57 <= _GEN_57;
    end
    if (reset) begin
      valids_58 <= 1'h0;
    end else if (io_branch) begin
      valids_58 <= _GEN_58;
    end
    if (reset) begin
      valids_59 <= 1'h0;
    end else if (io_branch) begin
      valids_59 <= _GEN_59;
    end
    if (reset) begin
      valids_60 <= 1'h0;
    end else if (io_branch) begin
      valids_60 <= _GEN_60;
    end
    if (reset) begin
      valids_61 <= 1'h0;
    end else if (io_branch) begin
      valids_61 <= _GEN_61;
    end
    if (reset) begin
      valids_62 <= 1'h0;
    end else if (io_branch) begin
      valids_62 <= _GEN_62;
    end
    if (reset) begin
      valids_63 <= 1'h0;
    end else if (io_branch) begin
      valids_63 <= _GEN_63;
    end
  end
endmodule
module BranchPredictor(
  input         clock,
  input         reset,
  input         io_branchInfo_branch,
  input         io_branchInfo_jump,
  input         io_branchInfo_taken,
  input  [4:0]  io_branchInfo_index,
  input  [31:0] io_branchInfo_pc,
  input  [31:0] io_branchInfo_target,
  input  [31:0] io_lookupPc,
  output        io_predTaken,
  output [31:0] io_predTarget,
  output [4:0]  io_predIndex
);
  wire  ghr_clock; // @[BranchPredictor.scala 21:19]
  wire  ghr_io_branch; // @[BranchPredictor.scala 21:19]
  wire  ghr_io_taken; // @[BranchPredictor.scala 21:19]
  wire [4:0] ghr_io_ghr; // @[BranchPredictor.scala 21:19]
  wire  pht_clock; // @[BranchPredictor.scala 22:19]
  wire  pht_reset; // @[BranchPredictor.scala 22:19]
  wire  pht_io_lastBranch; // @[BranchPredictor.scala 22:19]
  wire  pht_io_lastTaken; // @[BranchPredictor.scala 22:19]
  wire [4:0] pht_io_lastIndex; // @[BranchPredictor.scala 22:19]
  wire [4:0] pht_io_index; // @[BranchPredictor.scala 22:19]
  wire  pht_io_taken; // @[BranchPredictor.scala 22:19]
  wire  btb_clock; // @[BranchPredictor.scala 23:19]
  wire  btb_reset; // @[BranchPredictor.scala 23:19]
  wire  btb_io_branch; // @[BranchPredictor.scala 23:19]
  wire  btb_io_jump; // @[BranchPredictor.scala 23:19]
  wire [31:0] btb_io_pc; // @[BranchPredictor.scala 23:19]
  wire [31:0] btb_io_target; // @[BranchPredictor.scala 23:19]
  wire [31:0] btb_io_lookupPc; // @[BranchPredictor.scala 23:19]
  wire  btb_io_lookupBranch; // @[BranchPredictor.scala 23:19]
  wire  btb_io_lookupJump; // @[BranchPredictor.scala 23:19]
  wire [31:0] btb_io_lookupTarget; // @[BranchPredictor.scala 23:19]
  wire  _T_1 = pht_io_taken | btb_io_lookupJump; // @[BranchPredictor.scala 46:34]
  GHR ghr ( // @[BranchPredictor.scala 21:19]
    .clock(ghr_clock),
    .io_branch(ghr_io_branch),
    .io_taken(ghr_io_taken),
    .io_ghr(ghr_io_ghr)
  );
  PHT pht ( // @[BranchPredictor.scala 22:19]
    .clock(pht_clock),
    .reset(pht_reset),
    .io_lastBranch(pht_io_lastBranch),
    .io_lastTaken(pht_io_lastTaken),
    .io_lastIndex(pht_io_lastIndex),
    .io_index(pht_io_index),
    .io_taken(pht_io_taken)
  );
  BTB btb ( // @[BranchPredictor.scala 23:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_branch(btb_io_branch),
    .io_jump(btb_io_jump),
    .io_pc(btb_io_pc),
    .io_target(btb_io_target),
    .io_lookupPc(btb_io_lookupPc),
    .io_lookupBranch(btb_io_lookupBranch),
    .io_lookupJump(btb_io_lookupJump),
    .io_lookupTarget(btb_io_lookupTarget)
  );
  assign io_predTaken = btb_io_lookupBranch & _T_1; // @[BranchPredictor.scala 45:17]
  assign io_predTarget = btb_io_lookupTarget; // @[BranchPredictor.scala 47:17]
  assign io_predIndex = io_lookupPc[6:2] ^ ghr_io_ghr; // @[BranchPredictor.scala 48:17]
  assign ghr_clock = clock;
  assign ghr_io_branch = io_branchInfo_branch; // @[BranchPredictor.scala 26:17]
  assign ghr_io_taken = io_branchInfo_taken; // @[BranchPredictor.scala 27:17]
  assign pht_clock = clock;
  assign pht_reset = reset;
  assign pht_io_lastBranch = io_branchInfo_branch; // @[BranchPredictor.scala 32:21]
  assign pht_io_lastTaken = io_branchInfo_taken; // @[BranchPredictor.scala 33:21]
  assign pht_io_lastIndex = io_branchInfo_index; // @[BranchPredictor.scala 34:21]
  assign pht_io_index = io_lookupPc[6:2] ^ ghr_io_ghr; // @[BranchPredictor.scala 35:21]
  assign btb_clock = clock;
  assign btb_reset = reset;
  assign btb_io_branch = io_branchInfo_branch; // @[BranchPredictor.scala 38:19]
  assign btb_io_jump = io_branchInfo_jump; // @[BranchPredictor.scala 39:19]
  assign btb_io_pc = io_branchInfo_pc; // @[BranchPredictor.scala 40:19]
  assign btb_io_target = io_branchInfo_target; // @[BranchPredictor.scala 41:19]
  assign btb_io_lookupPc = io_lookupPc; // @[BranchPredictor.scala 42:19]
endmodule
module Fetch(
  input         clock,
  input         reset,
  input         io_flush,
  input         io_stall,
  output        io_stallReq,
  input  [31:0] io_flushPc,
  input         io_rom_valid,
  input         io_rom_fault,
  output [31:0] io_rom_addr,
  input         io_branch_branch,
  input         io_branch_jump,
  input         io_branch_taken,
  input  [4:0]  io_branch_index,
  input  [31:0] io_branch_pc,
  input  [31:0] io_branch_target,
  output        io_fetch_valid,
  output [31:0] io_fetch_pc,
  output        io_fetch_taken,
  output [31:0] io_fetch_target,
  output [4:0]  io_fetch_predIndex,
  output        io_fetch_pageFault
);
  wire  bpu_clock; // @[Fetch.scala 28:19]
  wire  bpu_reset; // @[Fetch.scala 28:19]
  wire  bpu_io_branchInfo_branch; // @[Fetch.scala 28:19]
  wire  bpu_io_branchInfo_jump; // @[Fetch.scala 28:19]
  wire  bpu_io_branchInfo_taken; // @[Fetch.scala 28:19]
  wire [4:0] bpu_io_branchInfo_index; // @[Fetch.scala 28:19]
  wire [31:0] bpu_io_branchInfo_pc; // @[Fetch.scala 28:19]
  wire [31:0] bpu_io_branchInfo_target; // @[Fetch.scala 28:19]
  wire [31:0] bpu_io_lookupPc; // @[Fetch.scala 28:19]
  wire  bpu_io_predTaken; // @[Fetch.scala 28:19]
  wire [31:0] bpu_io_predTarget; // @[Fetch.scala 28:19]
  wire [4:0] bpu_io_predIndex; // @[Fetch.scala 28:19]
  reg [31:0] pc; // @[Fetch.scala 25:19]
  reg [31:0] _RAND_0;
  wire [31:0] _T_1 = pc + 32'h4; // @[Fetch.scala 36:23]
  BranchPredictor bpu ( // @[Fetch.scala 28:19]
    .clock(bpu_clock),
    .reset(bpu_reset),
    .io_branchInfo_branch(bpu_io_branchInfo_branch),
    .io_branchInfo_jump(bpu_io_branchInfo_jump),
    .io_branchInfo_taken(bpu_io_branchInfo_taken),
    .io_branchInfo_index(bpu_io_branchInfo_index),
    .io_branchInfo_pc(bpu_io_branchInfo_pc),
    .io_branchInfo_target(bpu_io_branchInfo_target),
    .io_lookupPc(bpu_io_lookupPc),
    .io_predTaken(bpu_io_predTaken),
    .io_predTarget(bpu_io_predTarget),
    .io_predIndex(bpu_io_predIndex)
  );
  assign io_stallReq = ~io_rom_valid; // @[Fetch.scala 40:15]
  assign io_rom_addr = pc; // @[Fetch.scala 45:17]
  assign io_fetch_valid = io_rom_valid; // @[Fetch.scala 49:23]
  assign io_fetch_pc = pc; // @[Fetch.scala 50:23]
  assign io_fetch_taken = bpu_io_predTaken; // @[Fetch.scala 51:23]
  assign io_fetch_target = bpu_io_predTarget; // @[Fetch.scala 52:23]
  assign io_fetch_predIndex = bpu_io_predIndex; // @[Fetch.scala 53:23]
  assign io_fetch_pageFault = io_rom_fault; // @[Fetch.scala 54:23]
  assign bpu_clock = clock;
  assign bpu_reset = reset;
  assign bpu_io_branchInfo_branch = io_branch_branch; // @[Fetch.scala 29:21]
  assign bpu_io_branchInfo_jump = io_branch_jump; // @[Fetch.scala 29:21]
  assign bpu_io_branchInfo_taken = io_branch_taken; // @[Fetch.scala 29:21]
  assign bpu_io_branchInfo_index = io_branch_index; // @[Fetch.scala 29:21]
  assign bpu_io_branchInfo_pc = io_branch_pc; // @[Fetch.scala 29:21]
  assign bpu_io_branchInfo_target = io_branch_target; // @[Fetch.scala 29:21]
  assign bpu_io_lookupPc = pc; // @[Fetch.scala 30:21]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pc <= 32'h200;
    end else if (io_flush) begin
      pc <= io_flushPc;
    end else if (!(io_stall)) begin
      if (bpu_io_predTaken) begin
        pc <= bpu_io_predTarget;
      end else begin
        pc <= _T_1;
      end
    end
  end
endmodule
module MidStage(
  input         clock,
  input         reset,
  input         io_flush,
  input         io_stallPrev,
  input         io_stallNext,
  input         io_prev_valid,
  input  [31:0] io_prev_pc,
  input         io_prev_taken,
  input  [31:0] io_prev_target,
  input  [4:0]  io_prev_predIndex,
  input         io_prev_pageFault,
  output        io_next_valid,
  output [31:0] io_next_pc,
  output        io_next_taken,
  output [31:0] io_next_target,
  output [4:0]  io_next_predIndex,
  output        io_next_pageFault
);
  reg  ff_valid; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_0;
  reg [31:0] ff_pc; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_1;
  reg  ff_taken; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_2;
  reg [31:0] ff_target; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_3;
  reg [4:0] ff_predIndex; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_4;
  reg  ff_pageFault; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_5;
  wire  _T_1 = ~io_stallNext; // @[MidStage.scala 21:38]
  wire  _T_2 = io_stallPrev & _T_1; // @[MidStage.scala 21:35]
  wire  _T_3 = io_flush | _T_2; // @[MidStage.scala 21:18]
  wire  _T_5 = ~io_stallPrev; // @[MidStage.scala 23:15]
  assign io_next_valid = ff_valid; // @[MidStage.scala 27:11]
  assign io_next_pc = ff_pc; // @[MidStage.scala 27:11]
  assign io_next_taken = ff_taken; // @[MidStage.scala 27:11]
  assign io_next_target = ff_target; // @[MidStage.scala 27:11]
  assign io_next_predIndex = ff_predIndex; // @[MidStage.scala 27:11]
  assign io_next_pageFault = ff_pageFault; // @[MidStage.scala 27:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ff_pc = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ff_taken = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ff_target = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ff_predIndex = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ff_pageFault = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ff_valid <= 1'h0;
    end else if (_T_3) begin
      ff_valid <= 1'h0;
    end else if (_T_5) begin
      ff_valid <= io_prev_valid;
    end
    if (reset) begin
      ff_pc <= 32'h0;
    end else if (_T_3) begin
      ff_pc <= 32'h0;
    end else if (_T_5) begin
      ff_pc <= io_prev_pc;
    end
    if (reset) begin
      ff_taken <= 1'h0;
    end else if (_T_3) begin
      ff_taken <= 1'h0;
    end else if (_T_5) begin
      ff_taken <= io_prev_taken;
    end
    if (reset) begin
      ff_target <= 32'h0;
    end else if (_T_3) begin
      ff_target <= 32'h0;
    end else if (_T_5) begin
      ff_target <= io_prev_target;
    end
    if (reset) begin
      ff_predIndex <= 5'h0;
    end else if (_T_3) begin
      ff_predIndex <= 5'h0;
    end else if (_T_5) begin
      ff_predIndex <= io_prev_predIndex;
    end
    if (reset) begin
      ff_pageFault <= 1'h0;
    end else if (_T_3) begin
      ff_pageFault <= 1'h0;
    end else if (_T_5) begin
      ff_pageFault <= io_prev_pageFault;
    end
  end
endmodule
module Decoder(
  input         clock,
  input         io_fetch_valid,
  input  [31:0] io_fetch_pc,
  input         io_fetch_taken,
  input  [31:0] io_fetch_target,
  input  [4:0]  io_fetch_predIndex,
  input         io_fetch_pageFault,
  input  [31:0] io_inst,
  input         io_stallId,
  output        io_flushIf,
  output [31:0] io_flushPc,
  output        io_read1_en,
  output [4:0]  io_read1_addr,
  input  [31:0] io_read1_data,
  output        io_read2_en,
  output [4:0]  io_read2_addr,
  input  [31:0] io_read2_data,
  output        io_branch_branch,
  output        io_branch_jump,
  output        io_branch_taken,
  output [4:0]  io_branch_index,
  output [31:0] io_branch_pc,
  output [31:0] io_branch_target,
  output [3:0]  io_decoder_aluOp,
  output [31:0] io_decoder_opr1,
  output [31:0] io_decoder_opr2,
  output [3:0]  io_decoder_mduOp,
  output [4:0]  io_decoder_lsuOp,
  output [31:0] io_decoder_lsuData,
  output        io_decoder_regWen,
  output [4:0]  io_decoder_regWaddr,
  output [2:0]  io_decoder_csrOp,
  output [11:0] io_decoder_csrAddr,
  output [31:0] io_decoder_csrData,
  output [3:0]  io_decoder_excType,
  output [31:0] io_decoder_excValue,
  output        io_decoder_valid,
  output [31:0] io_decoder_inst,
  output [31:0] io_decoder_currentPc
);
  reg  stallDelay; // @[Decoder.scala 36:28]
  reg [31:0] _RAND_0;
  reg [31:0] lastInst; // @[Decoder.scala 37:24]
  reg [31:0] _RAND_1;
  wire  _T = ~io_fetch_valid; // @[Decoder.scala 38:25]
  wire [31:0] _T_1 = stallDelay ? lastInst : io_inst; // @[Decoder.scala 39:24]
  wire [31:0] inst = _T ? 32'h13 : _T_1; // @[Decoder.scala 38:24]
  wire  _T_2 = ~stallDelay; // @[Decoder.scala 40:9]
  wire [4:0] rd = inst[11:7]; // @[Decoder.scala 43:17]
  wire [4:0] rs1 = inst[19:15]; // @[Decoder.scala 44:17]
  wire [4:0] rs2 = inst[24:20]; // @[Decoder.scala 45:17]
  wire [31:0] _T_20 = inst & 32'hfe00707f; // @[Lookup.scala 31:38]
  wire  _T_21 = 32'h33 == _T_20; // @[Lookup.scala 31:38]
  wire [31:0] _T_22 = inst & 32'h707f; // @[Lookup.scala 31:38]
  wire  _T_23 = 32'h13 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_25 = 32'h40000033 == _T_20; // @[Lookup.scala 31:38]
  wire [31:0] _T_26 = inst & 32'h7f; // @[Lookup.scala 31:38]
  wire  _T_27 = 32'h37 == _T_26; // @[Lookup.scala 31:38]
  wire  _T_29 = 32'h17 == _T_26; // @[Lookup.scala 31:38]
  wire  _T_31 = 32'h4033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_33 = 32'h4013 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_35 = 32'h6033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_37 = 32'h6013 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_39 = 32'h7033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_41 = 32'h7013 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_43 = 32'h2033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_45 = 32'h2013 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_47 = 32'h3033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_49 = 32'h3013 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_51 = 32'h1033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_53 = 32'h1013 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_55 = 32'h5033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_57 = 32'h5013 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_59 = 32'h40005033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_61 = 32'h40005013 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_63 = 32'h63 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_65 = 32'h1063 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_67 = 32'h4063 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_69 = 32'h5063 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_71 = 32'h6063 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_73 = 32'h7063 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_75 = 32'h6f == _T_26; // @[Lookup.scala 31:38]
  wire  _T_77 = 32'h67 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_79 = 32'h3 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_81 = 32'h1003 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_83 = 32'h2003 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_85 = 32'h4003 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_87 = 32'h5003 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_89 = 32'h23 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_91 = 32'h1023 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_93 = 32'h2023 == _T_22; // @[Lookup.scala 31:38]
  wire [31:0] _T_94 = inst & 32'hf00fffff; // @[Lookup.scala 31:38]
  wire  _T_95 = 32'hf == _T_94; // @[Lookup.scala 31:38]
  wire  _T_97 = 32'h100f == inst; // @[Lookup.scala 31:38]
  wire  _T_99 = 32'h1073 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_101 = 32'h2073 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_103 = 32'h3073 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_105 = 32'h5073 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_107 = 32'h6073 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_109 = 32'h7073 == _T_22; // @[Lookup.scala 31:38]
  wire  _T_111 = 32'h2000033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_113 = 32'h2001033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_115 = 32'h2002033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_117 = 32'h2003033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_119 = 32'h2004033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_121 = 32'h2005033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_123 = 32'h2006033 == _T_20; // @[Lookup.scala 31:38]
  wire  _T_125 = 32'h2007033 == _T_20; // @[Lookup.scala 31:38]
  wire [31:0] _T_126 = inst & 32'hf9f0707f; // @[Lookup.scala 31:38]
  wire  _T_127 = 32'h1000202f == _T_126; // @[Lookup.scala 31:38]
  wire [31:0] _T_128 = inst & 32'hf800707f; // @[Lookup.scala 31:38]
  wire  _T_129 = 32'h1800202f == _T_128; // @[Lookup.scala 31:38]
  wire  _T_131 = 32'h800202f == _T_128; // @[Lookup.scala 31:38]
  wire  _T_133 = 32'h202f == _T_128; // @[Lookup.scala 31:38]
  wire  _T_135 = 32'h2000202f == _T_128; // @[Lookup.scala 31:38]
  wire  _T_137 = 32'h6000202f == _T_128; // @[Lookup.scala 31:38]
  wire  _T_139 = 32'h4000202f == _T_128; // @[Lookup.scala 31:38]
  wire  _T_141 = 32'h8000202f == _T_128; // @[Lookup.scala 31:38]
  wire  _T_143 = 32'ha000202f == _T_128; // @[Lookup.scala 31:38]
  wire  _T_145 = 32'hc000202f == _T_128; // @[Lookup.scala 31:38]
  wire  _T_147 = 32'he000202f == _T_128; // @[Lookup.scala 31:38]
  wire  _T_149 = 32'h73 == inst; // @[Lookup.scala 31:38]
  wire  _T_151 = 32'h100073 == inst; // @[Lookup.scala 31:38]
  wire  _T_153 = 32'h10200073 == inst; // @[Lookup.scala 31:38]
  wire  _T_155 = 32'h30200073 == inst; // @[Lookup.scala 31:38]
  wire  _T_157 = 32'h10500073 == inst; // @[Lookup.scala 31:38]
  wire [31:0] _T_158 = inst & 32'hfe007fff; // @[Lookup.scala 31:38]
  wire  _T_159 = 32'h12000073 == _T_158; // @[Lookup.scala 31:38]
  wire  _T_161 = _T_157 ? 1'h0 : _T_159; // @[Lookup.scala 33:37]
  wire  _T_162 = _T_155 ? 1'h0 : _T_161; // @[Lookup.scala 33:37]
  wire  _T_163 = _T_153 ? 1'h0 : _T_162; // @[Lookup.scala 33:37]
  wire  _T_164 = _T_151 ? 1'h0 : _T_163; // @[Lookup.scala 33:37]
  wire  _T_165 = _T_149 ? 1'h0 : _T_164; // @[Lookup.scala 33:37]
  wire  _T_166 = _T_147 | _T_165; // @[Lookup.scala 33:37]
  wire  _T_167 = _T_145 | _T_166; // @[Lookup.scala 33:37]
  wire  _T_168 = _T_143 | _T_167; // @[Lookup.scala 33:37]
  wire  _T_169 = _T_141 | _T_168; // @[Lookup.scala 33:37]
  wire  _T_170 = _T_139 | _T_169; // @[Lookup.scala 33:37]
  wire  _T_171 = _T_137 | _T_170; // @[Lookup.scala 33:37]
  wire  _T_172 = _T_135 | _T_171; // @[Lookup.scala 33:37]
  wire  _T_173 = _T_133 | _T_172; // @[Lookup.scala 33:37]
  wire  _T_174 = _T_131 | _T_173; // @[Lookup.scala 33:37]
  wire  _T_175 = _T_129 | _T_174; // @[Lookup.scala 33:37]
  wire  _T_176 = _T_127 | _T_175; // @[Lookup.scala 33:37]
  wire  _T_177 = _T_125 | _T_176; // @[Lookup.scala 33:37]
  wire  _T_178 = _T_123 | _T_177; // @[Lookup.scala 33:37]
  wire  _T_179 = _T_121 | _T_178; // @[Lookup.scala 33:37]
  wire  _T_180 = _T_119 | _T_179; // @[Lookup.scala 33:37]
  wire  _T_181 = _T_117 | _T_180; // @[Lookup.scala 33:37]
  wire  _T_182 = _T_115 | _T_181; // @[Lookup.scala 33:37]
  wire  _T_183 = _T_113 | _T_182; // @[Lookup.scala 33:37]
  wire  _T_184 = _T_111 | _T_183; // @[Lookup.scala 33:37]
  wire  _T_185 = _T_109 ? 1'h0 : _T_184; // @[Lookup.scala 33:37]
  wire  _T_186 = _T_107 ? 1'h0 : _T_185; // @[Lookup.scala 33:37]
  wire  _T_187 = _T_105 ? 1'h0 : _T_186; // @[Lookup.scala 33:37]
  wire  _T_188 = _T_103 | _T_187; // @[Lookup.scala 33:37]
  wire  _T_189 = _T_101 | _T_188; // @[Lookup.scala 33:37]
  wire  _T_190 = _T_99 | _T_189; // @[Lookup.scala 33:37]
  wire  _T_191 = _T_97 ? 1'h0 : _T_190; // @[Lookup.scala 33:37]
  wire  _T_192 = _T_95 ? 1'h0 : _T_191; // @[Lookup.scala 33:37]
  wire  _T_193 = _T_93 | _T_192; // @[Lookup.scala 33:37]
  wire  _T_194 = _T_91 | _T_193; // @[Lookup.scala 33:37]
  wire  _T_195 = _T_89 | _T_194; // @[Lookup.scala 33:37]
  wire  _T_196 = _T_87 | _T_195; // @[Lookup.scala 33:37]
  wire  _T_197 = _T_85 | _T_196; // @[Lookup.scala 33:37]
  wire  _T_198 = _T_83 | _T_197; // @[Lookup.scala 33:37]
  wire  _T_199 = _T_81 | _T_198; // @[Lookup.scala 33:37]
  wire  _T_200 = _T_79 | _T_199; // @[Lookup.scala 33:37]
  wire  _T_201 = _T_77 | _T_200; // @[Lookup.scala 33:37]
  wire  _T_202 = _T_75 ? 1'h0 : _T_201; // @[Lookup.scala 33:37]
  wire  _T_203 = _T_73 | _T_202; // @[Lookup.scala 33:37]
  wire  _T_204 = _T_71 | _T_203; // @[Lookup.scala 33:37]
  wire  _T_205 = _T_69 | _T_204; // @[Lookup.scala 33:37]
  wire  _T_206 = _T_67 | _T_205; // @[Lookup.scala 33:37]
  wire  _T_207 = _T_65 | _T_206; // @[Lookup.scala 33:37]
  wire  _T_208 = _T_63 | _T_207; // @[Lookup.scala 33:37]
  wire  _T_209 = _T_61 | _T_208; // @[Lookup.scala 33:37]
  wire  _T_210 = _T_59 | _T_209; // @[Lookup.scala 33:37]
  wire  _T_211 = _T_57 | _T_210; // @[Lookup.scala 33:37]
  wire  _T_212 = _T_55 | _T_211; // @[Lookup.scala 33:37]
  wire  _T_213 = _T_53 | _T_212; // @[Lookup.scala 33:37]
  wire  _T_214 = _T_51 | _T_213; // @[Lookup.scala 33:37]
  wire  _T_215 = _T_49 | _T_214; // @[Lookup.scala 33:37]
  wire  _T_216 = _T_47 | _T_215; // @[Lookup.scala 33:37]
  wire  _T_217 = _T_45 | _T_216; // @[Lookup.scala 33:37]
  wire  _T_218 = _T_43 | _T_217; // @[Lookup.scala 33:37]
  wire  _T_219 = _T_41 | _T_218; // @[Lookup.scala 33:37]
  wire  _T_220 = _T_39 | _T_219; // @[Lookup.scala 33:37]
  wire  _T_221 = _T_37 | _T_220; // @[Lookup.scala 33:37]
  wire  _T_222 = _T_35 | _T_221; // @[Lookup.scala 33:37]
  wire  _T_223 = _T_33 | _T_222; // @[Lookup.scala 33:37]
  wire  _T_224 = _T_31 | _T_223; // @[Lookup.scala 33:37]
  wire  _T_225 = _T_29 ? 1'h0 : _T_224; // @[Lookup.scala 33:37]
  wire  _T_226 = _T_27 ? 1'h0 : _T_225; // @[Lookup.scala 33:37]
  wire  _T_227 = _T_25 | _T_226; // @[Lookup.scala 33:37]
  wire  _T_228 = _T_23 | _T_227; // @[Lookup.scala 33:37]
  wire  regEn1 = _T_21 | _T_228; // @[Lookup.scala 33:37]
  wire  _T_245 = _T_127 ? 1'h0 : _T_175; // @[Lookup.scala 33:37]
  wire  _T_246 = _T_125 | _T_245; // @[Lookup.scala 33:37]
  wire  _T_247 = _T_123 | _T_246; // @[Lookup.scala 33:37]
  wire  _T_248 = _T_121 | _T_247; // @[Lookup.scala 33:37]
  wire  _T_249 = _T_119 | _T_248; // @[Lookup.scala 33:37]
  wire  _T_250 = _T_117 | _T_249; // @[Lookup.scala 33:37]
  wire  _T_251 = _T_115 | _T_250; // @[Lookup.scala 33:37]
  wire  _T_252 = _T_113 | _T_251; // @[Lookup.scala 33:37]
  wire  _T_253 = _T_111 | _T_252; // @[Lookup.scala 33:37]
  wire  _T_254 = _T_109 ? 1'h0 : _T_253; // @[Lookup.scala 33:37]
  wire  _T_255 = _T_107 ? 1'h0 : _T_254; // @[Lookup.scala 33:37]
  wire  _T_256 = _T_105 ? 1'h0 : _T_255; // @[Lookup.scala 33:37]
  wire  _T_257 = _T_103 ? 1'h0 : _T_256; // @[Lookup.scala 33:37]
  wire  _T_258 = _T_101 ? 1'h0 : _T_257; // @[Lookup.scala 33:37]
  wire  _T_259 = _T_99 ? 1'h0 : _T_258; // @[Lookup.scala 33:37]
  wire  _T_260 = _T_97 ? 1'h0 : _T_259; // @[Lookup.scala 33:37]
  wire  _T_261 = _T_95 ? 1'h0 : _T_260; // @[Lookup.scala 33:37]
  wire  _T_262 = _T_93 | _T_261; // @[Lookup.scala 33:37]
  wire  _T_263 = _T_91 | _T_262; // @[Lookup.scala 33:37]
  wire  _T_264 = _T_89 | _T_263; // @[Lookup.scala 33:37]
  wire  _T_265 = _T_87 ? 1'h0 : _T_264; // @[Lookup.scala 33:37]
  wire  _T_266 = _T_85 ? 1'h0 : _T_265; // @[Lookup.scala 33:37]
  wire  _T_267 = _T_83 ? 1'h0 : _T_266; // @[Lookup.scala 33:37]
  wire  _T_268 = _T_81 ? 1'h0 : _T_267; // @[Lookup.scala 33:37]
  wire  _T_269 = _T_79 ? 1'h0 : _T_268; // @[Lookup.scala 33:37]
  wire  _T_270 = _T_77 ? 1'h0 : _T_269; // @[Lookup.scala 33:37]
  wire  _T_271 = _T_75 ? 1'h0 : _T_270; // @[Lookup.scala 33:37]
  wire  _T_272 = _T_73 | _T_271; // @[Lookup.scala 33:37]
  wire  _T_273 = _T_71 | _T_272; // @[Lookup.scala 33:37]
  wire  _T_274 = _T_69 | _T_273; // @[Lookup.scala 33:37]
  wire  _T_275 = _T_67 | _T_274; // @[Lookup.scala 33:37]
  wire  _T_276 = _T_65 | _T_275; // @[Lookup.scala 33:37]
  wire  _T_277 = _T_63 | _T_276; // @[Lookup.scala 33:37]
  wire  _T_278 = _T_61 ? 1'h0 : _T_277; // @[Lookup.scala 33:37]
  wire  _T_279 = _T_59 | _T_278; // @[Lookup.scala 33:37]
  wire  _T_280 = _T_57 ? 1'h0 : _T_279; // @[Lookup.scala 33:37]
  wire  _T_281 = _T_55 | _T_280; // @[Lookup.scala 33:37]
  wire  _T_282 = _T_53 ? 1'h0 : _T_281; // @[Lookup.scala 33:37]
  wire  _T_283 = _T_51 | _T_282; // @[Lookup.scala 33:37]
  wire  _T_284 = _T_49 ? 1'h0 : _T_283; // @[Lookup.scala 33:37]
  wire  _T_285 = _T_47 | _T_284; // @[Lookup.scala 33:37]
  wire  _T_286 = _T_45 ? 1'h0 : _T_285; // @[Lookup.scala 33:37]
  wire  _T_287 = _T_43 | _T_286; // @[Lookup.scala 33:37]
  wire  _T_288 = _T_41 ? 1'h0 : _T_287; // @[Lookup.scala 33:37]
  wire  _T_289 = _T_39 | _T_288; // @[Lookup.scala 33:37]
  wire  _T_290 = _T_37 ? 1'h0 : _T_289; // @[Lookup.scala 33:37]
  wire  _T_291 = _T_35 | _T_290; // @[Lookup.scala 33:37]
  wire  _T_292 = _T_33 ? 1'h0 : _T_291; // @[Lookup.scala 33:37]
  wire  _T_293 = _T_31 | _T_292; // @[Lookup.scala 33:37]
  wire  _T_294 = _T_29 ? 1'h0 : _T_293; // @[Lookup.scala 33:37]
  wire  _T_295 = _T_27 ? 1'h0 : _T_294; // @[Lookup.scala 33:37]
  wire  _T_296 = _T_25 | _T_295; // @[Lookup.scala 33:37]
  wire  _T_297 = _T_23 ? 1'h0 : _T_296; // @[Lookup.scala 33:37]
  wire  _T_305 = _T_145 | _T_147; // @[Lookup.scala 33:37]
  wire  _T_306 = _T_143 | _T_305; // @[Lookup.scala 33:37]
  wire  _T_307 = _T_141 | _T_306; // @[Lookup.scala 33:37]
  wire  _T_308 = _T_139 | _T_307; // @[Lookup.scala 33:37]
  wire  _T_309 = _T_137 | _T_308; // @[Lookup.scala 33:37]
  wire  _T_310 = _T_135 | _T_309; // @[Lookup.scala 33:37]
  wire  _T_311 = _T_133 | _T_310; // @[Lookup.scala 33:37]
  wire  _T_312 = _T_131 | _T_311; // @[Lookup.scala 33:37]
  wire  _T_313 = _T_129 | _T_312; // @[Lookup.scala 33:37]
  wire  _T_314 = _T_127 | _T_313; // @[Lookup.scala 33:37]
  wire  _T_315 = _T_125 | _T_314; // @[Lookup.scala 33:37]
  wire  _T_316 = _T_123 | _T_315; // @[Lookup.scala 33:37]
  wire  _T_317 = _T_121 | _T_316; // @[Lookup.scala 33:37]
  wire  _T_318 = _T_119 | _T_317; // @[Lookup.scala 33:37]
  wire  _T_319 = _T_117 | _T_318; // @[Lookup.scala 33:37]
  wire  _T_320 = _T_115 | _T_319; // @[Lookup.scala 33:37]
  wire  _T_321 = _T_113 | _T_320; // @[Lookup.scala 33:37]
  wire  _T_322 = _T_111 | _T_321; // @[Lookup.scala 33:37]
  wire  _T_323 = _T_109 | _T_322; // @[Lookup.scala 33:37]
  wire  _T_324 = _T_107 | _T_323; // @[Lookup.scala 33:37]
  wire  _T_325 = _T_105 | _T_324; // @[Lookup.scala 33:37]
  wire  _T_326 = _T_103 | _T_325; // @[Lookup.scala 33:37]
  wire  _T_327 = _T_101 | _T_326; // @[Lookup.scala 33:37]
  wire  _T_328 = _T_99 | _T_327; // @[Lookup.scala 33:37]
  wire  _T_329 = _T_97 ? 1'h0 : _T_328; // @[Lookup.scala 33:37]
  wire  _T_330 = _T_95 ? 1'h0 : _T_329; // @[Lookup.scala 33:37]
  wire  _T_331 = _T_93 ? 1'h0 : _T_330; // @[Lookup.scala 33:37]
  wire  _T_332 = _T_91 ? 1'h0 : _T_331; // @[Lookup.scala 33:37]
  wire  _T_333 = _T_89 ? 1'h0 : _T_332; // @[Lookup.scala 33:37]
  wire  _T_334 = _T_87 | _T_333; // @[Lookup.scala 33:37]
  wire  _T_335 = _T_85 | _T_334; // @[Lookup.scala 33:37]
  wire  _T_336 = _T_83 | _T_335; // @[Lookup.scala 33:37]
  wire  _T_337 = _T_81 | _T_336; // @[Lookup.scala 33:37]
  wire  _T_338 = _T_79 | _T_337; // @[Lookup.scala 33:37]
  wire  _T_339 = _T_77 | _T_338; // @[Lookup.scala 33:37]
  wire  _T_340 = _T_75 | _T_339; // @[Lookup.scala 33:37]
  wire  _T_341 = _T_73 ? 1'h0 : _T_340; // @[Lookup.scala 33:37]
  wire  _T_342 = _T_71 ? 1'h0 : _T_341; // @[Lookup.scala 33:37]
  wire  _T_343 = _T_69 ? 1'h0 : _T_342; // @[Lookup.scala 33:37]
  wire  _T_344 = _T_67 ? 1'h0 : _T_343; // @[Lookup.scala 33:37]
  wire  _T_345 = _T_65 ? 1'h0 : _T_344; // @[Lookup.scala 33:37]
  wire  _T_346 = _T_63 ? 1'h0 : _T_345; // @[Lookup.scala 33:37]
  wire  _T_347 = _T_61 | _T_346; // @[Lookup.scala 33:37]
  wire  _T_348 = _T_59 | _T_347; // @[Lookup.scala 33:37]
  wire  _T_349 = _T_57 | _T_348; // @[Lookup.scala 33:37]
  wire  _T_350 = _T_55 | _T_349; // @[Lookup.scala 33:37]
  wire  _T_351 = _T_53 | _T_350; // @[Lookup.scala 33:37]
  wire  _T_352 = _T_51 | _T_351; // @[Lookup.scala 33:37]
  wire  _T_353 = _T_49 | _T_352; // @[Lookup.scala 33:37]
  wire  _T_354 = _T_47 | _T_353; // @[Lookup.scala 33:37]
  wire  _T_355 = _T_45 | _T_354; // @[Lookup.scala 33:37]
  wire  _T_356 = _T_43 | _T_355; // @[Lookup.scala 33:37]
  wire  _T_357 = _T_41 | _T_356; // @[Lookup.scala 33:37]
  wire  _T_358 = _T_39 | _T_357; // @[Lookup.scala 33:37]
  wire  _T_359 = _T_37 | _T_358; // @[Lookup.scala 33:37]
  wire  _T_360 = _T_35 | _T_359; // @[Lookup.scala 33:37]
  wire  _T_361 = _T_33 | _T_360; // @[Lookup.scala 33:37]
  wire  _T_362 = _T_31 | _T_361; // @[Lookup.scala 33:37]
  wire  _T_363 = _T_29 | _T_362; // @[Lookup.scala 33:37]
  wire  _T_364 = _T_27 | _T_363; // @[Lookup.scala 33:37]
  wire  _T_365 = _T_25 | _T_364; // @[Lookup.scala 33:37]
  wire  _T_366 = _T_23 | _T_365; // @[Lookup.scala 33:37]
  wire [3:0] _T_367 = _T_159 ? 4'h1 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_368 = _T_157 ? 4'h0 : _T_367; // @[Lookup.scala 33:37]
  wire [3:0] _T_369 = _T_155 ? 4'h0 : _T_368; // @[Lookup.scala 33:37]
  wire [3:0] _T_370 = _T_153 ? 4'h0 : _T_369; // @[Lookup.scala 33:37]
  wire [3:0] _T_371 = _T_151 ? 4'h0 : _T_370; // @[Lookup.scala 33:37]
  wire [3:0] _T_372 = _T_149 ? 4'h0 : _T_371; // @[Lookup.scala 33:37]
  wire [3:0] _T_373 = _T_147 ? 4'h1 : _T_372; // @[Lookup.scala 33:37]
  wire [3:0] _T_374 = _T_145 ? 4'h1 : _T_373; // @[Lookup.scala 33:37]
  wire [3:0] _T_375 = _T_143 ? 4'h1 : _T_374; // @[Lookup.scala 33:37]
  wire [3:0] _T_376 = _T_141 ? 4'h1 : _T_375; // @[Lookup.scala 33:37]
  wire [3:0] _T_377 = _T_139 ? 4'h1 : _T_376; // @[Lookup.scala 33:37]
  wire [3:0] _T_378 = _T_137 ? 4'h1 : _T_377; // @[Lookup.scala 33:37]
  wire [3:0] _T_379 = _T_135 ? 4'h1 : _T_378; // @[Lookup.scala 33:37]
  wire [3:0] _T_380 = _T_133 ? 4'h1 : _T_379; // @[Lookup.scala 33:37]
  wire [3:0] _T_381 = _T_131 ? 4'h1 : _T_380; // @[Lookup.scala 33:37]
  wire [3:0] _T_382 = _T_129 ? 4'h1 : _T_381; // @[Lookup.scala 33:37]
  wire [3:0] _T_383 = _T_127 ? 4'h1 : _T_382; // @[Lookup.scala 33:37]
  wire [3:0] _T_384 = _T_125 ? 4'h1 : _T_383; // @[Lookup.scala 33:37]
  wire [3:0] _T_385 = _T_123 ? 4'h1 : _T_384; // @[Lookup.scala 33:37]
  wire [3:0] _T_386 = _T_121 ? 4'h1 : _T_385; // @[Lookup.scala 33:37]
  wire [3:0] _T_387 = _T_119 ? 4'h1 : _T_386; // @[Lookup.scala 33:37]
  wire [3:0] _T_388 = _T_117 ? 4'h1 : _T_387; // @[Lookup.scala 33:37]
  wire [3:0] _T_389 = _T_115 ? 4'h1 : _T_388; // @[Lookup.scala 33:37]
  wire [3:0] _T_390 = _T_113 ? 4'h1 : _T_389; // @[Lookup.scala 33:37]
  wire [3:0] _T_391 = _T_111 ? 4'h1 : _T_390; // @[Lookup.scala 33:37]
  wire [3:0] _T_392 = _T_109 ? 4'h0 : _T_391; // @[Lookup.scala 33:37]
  wire [3:0] _T_393 = _T_107 ? 4'h0 : _T_392; // @[Lookup.scala 33:37]
  wire [3:0] _T_394 = _T_105 ? 4'h0 : _T_393; // @[Lookup.scala 33:37]
  wire [3:0] _T_395 = _T_103 ? 4'h0 : _T_394; // @[Lookup.scala 33:37]
  wire [3:0] _T_396 = _T_101 ? 4'h0 : _T_395; // @[Lookup.scala 33:37]
  wire [3:0] _T_397 = _T_99 ? 4'h0 : _T_396; // @[Lookup.scala 33:37]
  wire [3:0] _T_398 = _T_97 ? 4'h0 : _T_397; // @[Lookup.scala 33:37]
  wire [3:0] _T_399 = _T_95 ? 4'h0 : _T_398; // @[Lookup.scala 33:37]
  wire [3:0] _T_400 = _T_93 ? 4'h1 : _T_399; // @[Lookup.scala 33:37]
  wire [3:0] _T_401 = _T_91 ? 4'h1 : _T_400; // @[Lookup.scala 33:37]
  wire [3:0] _T_402 = _T_89 ? 4'h1 : _T_401; // @[Lookup.scala 33:37]
  wire [3:0] _T_403 = _T_87 ? 4'h1 : _T_402; // @[Lookup.scala 33:37]
  wire [3:0] _T_404 = _T_85 ? 4'h1 : _T_403; // @[Lookup.scala 33:37]
  wire [3:0] _T_405 = _T_83 ? 4'h1 : _T_404; // @[Lookup.scala 33:37]
  wire [3:0] _T_406 = _T_81 ? 4'h1 : _T_405; // @[Lookup.scala 33:37]
  wire [3:0] _T_407 = _T_79 ? 4'h1 : _T_406; // @[Lookup.scala 33:37]
  wire [3:0] _T_408 = _T_77 ? 4'h7 : _T_407; // @[Lookup.scala 33:37]
  wire [3:0] _T_409 = _T_75 ? 4'h7 : _T_408; // @[Lookup.scala 33:37]
  wire [3:0] _T_410 = _T_73 ? 4'h0 : _T_409; // @[Lookup.scala 33:37]
  wire [3:0] _T_411 = _T_71 ? 4'h0 : _T_410; // @[Lookup.scala 33:37]
  wire [3:0] _T_412 = _T_69 ? 4'h0 : _T_411; // @[Lookup.scala 33:37]
  wire [3:0] _T_413 = _T_67 ? 4'h0 : _T_412; // @[Lookup.scala 33:37]
  wire [3:0] _T_414 = _T_65 ? 4'h0 : _T_413; // @[Lookup.scala 33:37]
  wire [3:0] _T_415 = _T_63 ? 4'h0 : _T_414; // @[Lookup.scala 33:37]
  wire [3:0] _T_416 = _T_61 ? 4'h1 : _T_415; // @[Lookup.scala 33:37]
  wire [3:0] _T_417 = _T_59 ? 4'h1 : _T_416; // @[Lookup.scala 33:37]
  wire [3:0] _T_418 = _T_57 ? 4'h1 : _T_417; // @[Lookup.scala 33:37]
  wire [3:0] _T_419 = _T_55 ? 4'h1 : _T_418; // @[Lookup.scala 33:37]
  wire [3:0] _T_420 = _T_53 ? 4'h1 : _T_419; // @[Lookup.scala 33:37]
  wire [3:0] _T_421 = _T_51 ? 4'h1 : _T_420; // @[Lookup.scala 33:37]
  wire [3:0] _T_422 = _T_49 ? 4'h1 : _T_421; // @[Lookup.scala 33:37]
  wire [3:0] _T_423 = _T_47 ? 4'h1 : _T_422; // @[Lookup.scala 33:37]
  wire [3:0] _T_424 = _T_45 ? 4'h1 : _T_423; // @[Lookup.scala 33:37]
  wire [3:0] _T_425 = _T_43 ? 4'h1 : _T_424; // @[Lookup.scala 33:37]
  wire [3:0] _T_426 = _T_41 ? 4'h1 : _T_425; // @[Lookup.scala 33:37]
  wire [3:0] _T_427 = _T_39 ? 4'h1 : _T_426; // @[Lookup.scala 33:37]
  wire [3:0] _T_428 = _T_37 ? 4'h1 : _T_427; // @[Lookup.scala 33:37]
  wire [3:0] _T_429 = _T_35 ? 4'h1 : _T_428; // @[Lookup.scala 33:37]
  wire [3:0] _T_430 = _T_33 ? 4'h1 : _T_429; // @[Lookup.scala 33:37]
  wire [3:0] _T_431 = _T_31 ? 4'h1 : _T_430; // @[Lookup.scala 33:37]
  wire [3:0] _T_432 = _T_29 ? 4'h7 : _T_431; // @[Lookup.scala 33:37]
  wire [3:0] _T_433 = _T_27 ? 4'h0 : _T_432; // @[Lookup.scala 33:37]
  wire [3:0] _T_434 = _T_25 ? 4'h1 : _T_433; // @[Lookup.scala 33:37]
  wire [3:0] _T_435 = _T_23 ? 4'h1 : _T_434; // @[Lookup.scala 33:37]
  wire [3:0] aluSrc1 = _T_21 ? 4'h1 : _T_435; // @[Lookup.scala 33:37]
  wire [3:0] _T_453 = _T_125 ? 4'h2 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_454 = _T_123 ? 4'h2 : _T_453; // @[Lookup.scala 33:37]
  wire [3:0] _T_455 = _T_121 ? 4'h2 : _T_454; // @[Lookup.scala 33:37]
  wire [3:0] _T_456 = _T_119 ? 4'h2 : _T_455; // @[Lookup.scala 33:37]
  wire [3:0] _T_457 = _T_117 ? 4'h2 : _T_456; // @[Lookup.scala 33:37]
  wire [3:0] _T_458 = _T_115 ? 4'h2 : _T_457; // @[Lookup.scala 33:37]
  wire [3:0] _T_459 = _T_113 ? 4'h2 : _T_458; // @[Lookup.scala 33:37]
  wire [3:0] _T_460 = _T_111 ? 4'h2 : _T_459; // @[Lookup.scala 33:37]
  wire [3:0] _T_461 = _T_109 ? 4'h0 : _T_460; // @[Lookup.scala 33:37]
  wire [3:0] _T_462 = _T_107 ? 4'h0 : _T_461; // @[Lookup.scala 33:37]
  wire [3:0] _T_463 = _T_105 ? 4'h0 : _T_462; // @[Lookup.scala 33:37]
  wire [3:0] _T_464 = _T_103 ? 4'h0 : _T_463; // @[Lookup.scala 33:37]
  wire [3:0] _T_465 = _T_101 ? 4'h0 : _T_464; // @[Lookup.scala 33:37]
  wire [3:0] _T_466 = _T_99 ? 4'h0 : _T_465; // @[Lookup.scala 33:37]
  wire [3:0] _T_467 = _T_97 ? 4'h0 : _T_466; // @[Lookup.scala 33:37]
  wire [3:0] _T_468 = _T_95 ? 4'h3 : _T_467; // @[Lookup.scala 33:37]
  wire [3:0] _T_469 = _T_93 ? 4'h4 : _T_468; // @[Lookup.scala 33:37]
  wire [3:0] _T_470 = _T_91 ? 4'h4 : _T_469; // @[Lookup.scala 33:37]
  wire [3:0] _T_471 = _T_89 ? 4'h4 : _T_470; // @[Lookup.scala 33:37]
  wire [3:0] _T_472 = _T_87 ? 4'h3 : _T_471; // @[Lookup.scala 33:37]
  wire [3:0] _T_473 = _T_85 ? 4'h3 : _T_472; // @[Lookup.scala 33:37]
  wire [3:0] _T_474 = _T_83 ? 4'h3 : _T_473; // @[Lookup.scala 33:37]
  wire [3:0] _T_475 = _T_81 ? 4'h3 : _T_474; // @[Lookup.scala 33:37]
  wire [3:0] _T_476 = _T_79 ? 4'h3 : _T_475; // @[Lookup.scala 33:37]
  wire [3:0] _T_477 = _T_77 ? 4'h8 : _T_476; // @[Lookup.scala 33:37]
  wire [3:0] _T_478 = _T_75 ? 4'h8 : _T_477; // @[Lookup.scala 33:37]
  wire [3:0] _T_479 = _T_73 ? 4'h0 : _T_478; // @[Lookup.scala 33:37]
  wire [3:0] _T_480 = _T_71 ? 4'h0 : _T_479; // @[Lookup.scala 33:37]
  wire [3:0] _T_481 = _T_69 ? 4'h0 : _T_480; // @[Lookup.scala 33:37]
  wire [3:0] _T_482 = _T_67 ? 4'h0 : _T_481; // @[Lookup.scala 33:37]
  wire [3:0] _T_483 = _T_65 ? 4'h0 : _T_482; // @[Lookup.scala 33:37]
  wire [3:0] _T_484 = _T_63 ? 4'h0 : _T_483; // @[Lookup.scala 33:37]
  wire [3:0] _T_485 = _T_61 ? 4'h6 : _T_484; // @[Lookup.scala 33:37]
  wire [3:0] _T_486 = _T_59 ? 4'h2 : _T_485; // @[Lookup.scala 33:37]
  wire [3:0] _T_487 = _T_57 ? 4'h6 : _T_486; // @[Lookup.scala 33:37]
  wire [3:0] _T_488 = _T_55 ? 4'h2 : _T_487; // @[Lookup.scala 33:37]
  wire [3:0] _T_489 = _T_53 ? 4'h6 : _T_488; // @[Lookup.scala 33:37]
  wire [3:0] _T_490 = _T_51 ? 4'h2 : _T_489; // @[Lookup.scala 33:37]
  wire [3:0] _T_491 = _T_49 ? 4'h3 : _T_490; // @[Lookup.scala 33:37]
  wire [3:0] _T_492 = _T_47 ? 4'h2 : _T_491; // @[Lookup.scala 33:37]
  wire [3:0] _T_493 = _T_45 ? 4'h3 : _T_492; // @[Lookup.scala 33:37]
  wire [3:0] _T_494 = _T_43 ? 4'h2 : _T_493; // @[Lookup.scala 33:37]
  wire [3:0] _T_495 = _T_41 ? 4'h3 : _T_494; // @[Lookup.scala 33:37]
  wire [3:0] _T_496 = _T_39 ? 4'h2 : _T_495; // @[Lookup.scala 33:37]
  wire [3:0] _T_497 = _T_37 ? 4'h3 : _T_496; // @[Lookup.scala 33:37]
  wire [3:0] _T_498 = _T_35 ? 4'h2 : _T_497; // @[Lookup.scala 33:37]
  wire [3:0] _T_499 = _T_33 ? 4'h3 : _T_498; // @[Lookup.scala 33:37]
  wire [3:0] _T_500 = _T_31 ? 4'h2 : _T_499; // @[Lookup.scala 33:37]
  wire [3:0] _T_501 = _T_29 ? 4'h5 : _T_500; // @[Lookup.scala 33:37]
  wire [3:0] _T_502 = _T_27 ? 4'h5 : _T_501; // @[Lookup.scala 33:37]
  wire [3:0] _T_503 = _T_25 ? 4'h2 : _T_502; // @[Lookup.scala 33:37]
  wire [3:0] _T_504 = _T_23 ? 4'h3 : _T_503; // @[Lookup.scala 33:37]
  wire [3:0] aluSrc2 = _T_21 ? 4'h2 : _T_504; // @[Lookup.scala 33:37]
  wire [3:0] _T_505 = _T_159 ? 4'h3 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_506 = _T_157 ? 4'h0 : _T_505; // @[Lookup.scala 33:37]
  wire [3:0] _T_507 = _T_155 ? 4'h0 : _T_506; // @[Lookup.scala 33:37]
  wire [3:0] _T_508 = _T_153 ? 4'h0 : _T_507; // @[Lookup.scala 33:37]
  wire [3:0] _T_509 = _T_151 ? 4'h0 : _T_508; // @[Lookup.scala 33:37]
  wire [3:0] _T_510 = _T_149 ? 4'h0 : _T_509; // @[Lookup.scala 33:37]
  wire [3:0] _T_511 = _T_147 ? 4'h3 : _T_510; // @[Lookup.scala 33:37]
  wire [3:0] _T_512 = _T_145 ? 4'h3 : _T_511; // @[Lookup.scala 33:37]
  wire [3:0] _T_513 = _T_143 ? 4'h3 : _T_512; // @[Lookup.scala 33:37]
  wire [3:0] _T_514 = _T_141 ? 4'h3 : _T_513; // @[Lookup.scala 33:37]
  wire [3:0] _T_515 = _T_139 ? 4'h3 : _T_514; // @[Lookup.scala 33:37]
  wire [3:0] _T_516 = _T_137 ? 4'h3 : _T_515; // @[Lookup.scala 33:37]
  wire [3:0] _T_517 = _T_135 ? 4'h3 : _T_516; // @[Lookup.scala 33:37]
  wire [3:0] _T_518 = _T_133 ? 4'h3 : _T_517; // @[Lookup.scala 33:37]
  wire [3:0] _T_519 = _T_131 ? 4'h3 : _T_518; // @[Lookup.scala 33:37]
  wire [3:0] _T_520 = _T_129 ? 4'h3 : _T_519; // @[Lookup.scala 33:37]
  wire [3:0] _T_521 = _T_127 ? 4'h3 : _T_520; // @[Lookup.scala 33:37]
  wire [3:0] _T_522 = _T_125 ? 4'h0 : _T_521; // @[Lookup.scala 33:37]
  wire [3:0] _T_523 = _T_123 ? 4'h0 : _T_522; // @[Lookup.scala 33:37]
  wire [3:0] _T_524 = _T_121 ? 4'h0 : _T_523; // @[Lookup.scala 33:37]
  wire [3:0] _T_525 = _T_119 ? 4'h0 : _T_524; // @[Lookup.scala 33:37]
  wire [3:0] _T_526 = _T_117 ? 4'h0 : _T_525; // @[Lookup.scala 33:37]
  wire [3:0] _T_527 = _T_115 ? 4'h0 : _T_526; // @[Lookup.scala 33:37]
  wire [3:0] _T_528 = _T_113 ? 4'h0 : _T_527; // @[Lookup.scala 33:37]
  wire [3:0] _T_529 = _T_111 ? 4'h0 : _T_528; // @[Lookup.scala 33:37]
  wire [3:0] _T_530 = _T_109 ? 4'h0 : _T_529; // @[Lookup.scala 33:37]
  wire [3:0] _T_531 = _T_107 ? 4'h0 : _T_530; // @[Lookup.scala 33:37]
  wire [3:0] _T_532 = _T_105 ? 4'h0 : _T_531; // @[Lookup.scala 33:37]
  wire [3:0] _T_533 = _T_103 ? 4'h0 : _T_532; // @[Lookup.scala 33:37]
  wire [3:0] _T_534 = _T_101 ? 4'h0 : _T_533; // @[Lookup.scala 33:37]
  wire [3:0] _T_535 = _T_99 ? 4'h0 : _T_534; // @[Lookup.scala 33:37]
  wire [3:0] _T_536 = _T_97 ? 4'h0 : _T_535; // @[Lookup.scala 33:37]
  wire [3:0] _T_537 = _T_95 ? 4'h3 : _T_536; // @[Lookup.scala 33:37]
  wire [3:0] _T_538 = _T_93 ? 4'h0 : _T_537; // @[Lookup.scala 33:37]
  wire [3:0] _T_539 = _T_91 ? 4'h0 : _T_538; // @[Lookup.scala 33:37]
  wire [3:0] _T_540 = _T_89 ? 4'h0 : _T_539; // @[Lookup.scala 33:37]
  wire [3:0] _T_541 = _T_87 ? 4'h0 : _T_540; // @[Lookup.scala 33:37]
  wire [3:0] _T_542 = _T_85 ? 4'h0 : _T_541; // @[Lookup.scala 33:37]
  wire [3:0] _T_543 = _T_83 ? 4'h0 : _T_542; // @[Lookup.scala 33:37]
  wire [3:0] _T_544 = _T_81 ? 4'h0 : _T_543; // @[Lookup.scala 33:37]
  wire [3:0] _T_545 = _T_79 ? 4'h0 : _T_544; // @[Lookup.scala 33:37]
  wire [3:0] _T_546 = _T_77 ? 4'h0 : _T_545; // @[Lookup.scala 33:37]
  wire [3:0] _T_547 = _T_75 ? 4'h0 : _T_546; // @[Lookup.scala 33:37]
  wire [3:0] _T_548 = _T_73 ? 4'h0 : _T_547; // @[Lookup.scala 33:37]
  wire [3:0] _T_549 = _T_71 ? 4'h0 : _T_548; // @[Lookup.scala 33:37]
  wire [3:0] _T_550 = _T_69 ? 4'h0 : _T_549; // @[Lookup.scala 33:37]
  wire [3:0] _T_551 = _T_67 ? 4'h0 : _T_550; // @[Lookup.scala 33:37]
  wire [3:0] _T_552 = _T_65 ? 4'h0 : _T_551; // @[Lookup.scala 33:37]
  wire [3:0] _T_553 = _T_63 ? 4'h0 : _T_552; // @[Lookup.scala 33:37]
  wire [3:0] _T_554 = _T_61 ? 4'h9 : _T_553; // @[Lookup.scala 33:37]
  wire [3:0] _T_555 = _T_59 ? 4'h9 : _T_554; // @[Lookup.scala 33:37]
  wire [3:0] _T_556 = _T_57 ? 4'h8 : _T_555; // @[Lookup.scala 33:37]
  wire [3:0] _T_557 = _T_55 ? 4'h8 : _T_556; // @[Lookup.scala 33:37]
  wire [3:0] _T_558 = _T_53 ? 4'h7 : _T_557; // @[Lookup.scala 33:37]
  wire [3:0] _T_559 = _T_51 ? 4'h7 : _T_558; // @[Lookup.scala 33:37]
  wire [3:0] _T_560 = _T_49 ? 4'h6 : _T_559; // @[Lookup.scala 33:37]
  wire [3:0] _T_561 = _T_47 ? 4'h6 : _T_560; // @[Lookup.scala 33:37]
  wire [3:0] _T_562 = _T_45 ? 4'h5 : _T_561; // @[Lookup.scala 33:37]
  wire [3:0] _T_563 = _T_43 ? 4'h5 : _T_562; // @[Lookup.scala 33:37]
  wire [3:0] _T_564 = _T_41 ? 4'h4 : _T_563; // @[Lookup.scala 33:37]
  wire [3:0] _T_565 = _T_39 ? 4'h4 : _T_564; // @[Lookup.scala 33:37]
  wire [3:0] _T_566 = _T_37 ? 4'h3 : _T_565; // @[Lookup.scala 33:37]
  wire [3:0] _T_567 = _T_35 ? 4'h3 : _T_566; // @[Lookup.scala 33:37]
  wire [3:0] _T_568 = _T_33 ? 4'h2 : _T_567; // @[Lookup.scala 33:37]
  wire [3:0] _T_569 = _T_31 ? 4'h2 : _T_568; // @[Lookup.scala 33:37]
  wire [3:0] _T_570 = _T_29 ? 4'h0 : _T_569; // @[Lookup.scala 33:37]
  wire [3:0] _T_571 = _T_27 ? 4'h3 : _T_570; // @[Lookup.scala 33:37]
  wire [3:0] _T_572 = _T_25 ? 4'h1 : _T_571; // @[Lookup.scala 33:37]
  wire [3:0] _T_573 = _T_23 ? 4'h0 : _T_572; // @[Lookup.scala 33:37]
  wire [2:0] _T_615 = _T_77 ? 3'h1 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_616 = _T_75 ? 3'h1 : _T_615; // @[Lookup.scala 33:37]
  wire [2:0] _T_617 = _T_73 ? 3'h7 : _T_616; // @[Lookup.scala 33:37]
  wire [2:0] _T_618 = _T_71 ? 3'h6 : _T_617; // @[Lookup.scala 33:37]
  wire [2:0] _T_619 = _T_69 ? 3'h5 : _T_618; // @[Lookup.scala 33:37]
  wire [2:0] _T_620 = _T_67 ? 3'h4 : _T_619; // @[Lookup.scala 33:37]
  wire [2:0] _T_621 = _T_65 ? 3'h3 : _T_620; // @[Lookup.scala 33:37]
  wire [2:0] _T_622 = _T_63 ? 3'h2 : _T_621; // @[Lookup.scala 33:37]
  wire [2:0] _T_623 = _T_61 ? 3'h0 : _T_622; // @[Lookup.scala 33:37]
  wire [2:0] _T_624 = _T_59 ? 3'h0 : _T_623; // @[Lookup.scala 33:37]
  wire [2:0] _T_625 = _T_57 ? 3'h0 : _T_624; // @[Lookup.scala 33:37]
  wire [2:0] _T_626 = _T_55 ? 3'h0 : _T_625; // @[Lookup.scala 33:37]
  wire [2:0] _T_627 = _T_53 ? 3'h0 : _T_626; // @[Lookup.scala 33:37]
  wire [2:0] _T_628 = _T_51 ? 3'h0 : _T_627; // @[Lookup.scala 33:37]
  wire [2:0] _T_629 = _T_49 ? 3'h0 : _T_628; // @[Lookup.scala 33:37]
  wire [2:0] _T_630 = _T_47 ? 3'h0 : _T_629; // @[Lookup.scala 33:37]
  wire [2:0] _T_631 = _T_45 ? 3'h0 : _T_630; // @[Lookup.scala 33:37]
  wire [2:0] _T_632 = _T_43 ? 3'h0 : _T_631; // @[Lookup.scala 33:37]
  wire [2:0] _T_633 = _T_41 ? 3'h0 : _T_632; // @[Lookup.scala 33:37]
  wire [2:0] _T_634 = _T_39 ? 3'h0 : _T_633; // @[Lookup.scala 33:37]
  wire [2:0] _T_635 = _T_37 ? 3'h0 : _T_634; // @[Lookup.scala 33:37]
  wire [2:0] _T_636 = _T_35 ? 3'h0 : _T_635; // @[Lookup.scala 33:37]
  wire [2:0] _T_637 = _T_33 ? 3'h0 : _T_636; // @[Lookup.scala 33:37]
  wire [2:0] _T_638 = _T_31 ? 3'h0 : _T_637; // @[Lookup.scala 33:37]
  wire [2:0] _T_639 = _T_29 ? 3'h0 : _T_638; // @[Lookup.scala 33:37]
  wire [2:0] _T_640 = _T_27 ? 3'h0 : _T_639; // @[Lookup.scala 33:37]
  wire [2:0] _T_641 = _T_25 ? 3'h0 : _T_640; // @[Lookup.scala 33:37]
  wire [2:0] _T_642 = _T_23 ? 3'h0 : _T_641; // @[Lookup.scala 33:37]
  wire [2:0] branchFlag = _T_21 ? 3'h0 : _T_642; // @[Lookup.scala 33:37]
  wire [4:0] _T_643 = _T_159 ? 5'h16 : 5'h0; // @[Lookup.scala 33:37]
  wire [4:0] _T_644 = _T_157 ? 5'h0 : _T_643; // @[Lookup.scala 33:37]
  wire [4:0] _T_645 = _T_155 ? 5'h0 : _T_644; // @[Lookup.scala 33:37]
  wire [4:0] _T_646 = _T_153 ? 5'h0 : _T_645; // @[Lookup.scala 33:37]
  wire [4:0] _T_647 = _T_151 ? 5'h0 : _T_646; // @[Lookup.scala 33:37]
  wire [4:0] _T_648 = _T_149 ? 5'h0 : _T_647; // @[Lookup.scala 33:37]
  wire [4:0] _T_649 = _T_147 ? 5'h13 : _T_648; // @[Lookup.scala 33:37]
  wire [4:0] _T_650 = _T_145 ? 5'h12 : _T_649; // @[Lookup.scala 33:37]
  wire [4:0] _T_651 = _T_143 ? 5'h11 : _T_650; // @[Lookup.scala 33:37]
  wire [4:0] _T_652 = _T_141 ? 5'h10 : _T_651; // @[Lookup.scala 33:37]
  wire [4:0] _T_653 = _T_139 ? 5'hf : _T_652; // @[Lookup.scala 33:37]
  wire [4:0] _T_654 = _T_137 ? 5'he : _T_653; // @[Lookup.scala 33:37]
  wire [4:0] _T_655 = _T_135 ? 5'hd : _T_654; // @[Lookup.scala 33:37]
  wire [4:0] _T_656 = _T_133 ? 5'hc : _T_655; // @[Lookup.scala 33:37]
  wire [4:0] _T_657 = _T_131 ? 5'hb : _T_656; // @[Lookup.scala 33:37]
  wire [4:0] _T_658 = _T_129 ? 5'ha : _T_657; // @[Lookup.scala 33:37]
  wire [4:0] _T_659 = _T_127 ? 5'h9 : _T_658; // @[Lookup.scala 33:37]
  wire [4:0] _T_660 = _T_125 ? 5'h0 : _T_659; // @[Lookup.scala 33:37]
  wire [4:0] _T_661 = _T_123 ? 5'h0 : _T_660; // @[Lookup.scala 33:37]
  wire [4:0] _T_662 = _T_121 ? 5'h0 : _T_661; // @[Lookup.scala 33:37]
  wire [4:0] _T_663 = _T_119 ? 5'h0 : _T_662; // @[Lookup.scala 33:37]
  wire [4:0] _T_664 = _T_117 ? 5'h0 : _T_663; // @[Lookup.scala 33:37]
  wire [4:0] _T_665 = _T_115 ? 5'h0 : _T_664; // @[Lookup.scala 33:37]
  wire [4:0] _T_666 = _T_113 ? 5'h0 : _T_665; // @[Lookup.scala 33:37]
  wire [4:0] _T_667 = _T_111 ? 5'h0 : _T_666; // @[Lookup.scala 33:37]
  wire [4:0] _T_668 = _T_109 ? 5'h0 : _T_667; // @[Lookup.scala 33:37]
  wire [4:0] _T_669 = _T_107 ? 5'h0 : _T_668; // @[Lookup.scala 33:37]
  wire [4:0] _T_670 = _T_105 ? 5'h0 : _T_669; // @[Lookup.scala 33:37]
  wire [4:0] _T_671 = _T_103 ? 5'h0 : _T_670; // @[Lookup.scala 33:37]
  wire [4:0] _T_672 = _T_101 ? 5'h0 : _T_671; // @[Lookup.scala 33:37]
  wire [4:0] _T_673 = _T_99 ? 5'h0 : _T_672; // @[Lookup.scala 33:37]
  wire [4:0] _T_674 = _T_97 ? 5'h15 : _T_673; // @[Lookup.scala 33:37]
  wire [4:0] _T_675 = _T_95 ? 5'h14 : _T_674; // @[Lookup.scala 33:37]
  wire [4:0] _T_676 = _T_93 ? 5'h8 : _T_675; // @[Lookup.scala 33:37]
  wire [4:0] _T_677 = _T_91 ? 5'h7 : _T_676; // @[Lookup.scala 33:37]
  wire [4:0] _T_678 = _T_89 ? 5'h6 : _T_677; // @[Lookup.scala 33:37]
  wire [4:0] _T_679 = _T_87 ? 5'h5 : _T_678; // @[Lookup.scala 33:37]
  wire [4:0] _T_680 = _T_85 ? 5'h4 : _T_679; // @[Lookup.scala 33:37]
  wire [4:0] _T_681 = _T_83 ? 5'h3 : _T_680; // @[Lookup.scala 33:37]
  wire [4:0] _T_682 = _T_81 ? 5'h2 : _T_681; // @[Lookup.scala 33:37]
  wire [4:0] _T_683 = _T_79 ? 5'h1 : _T_682; // @[Lookup.scala 33:37]
  wire [4:0] _T_684 = _T_77 ? 5'h0 : _T_683; // @[Lookup.scala 33:37]
  wire [4:0] _T_685 = _T_75 ? 5'h0 : _T_684; // @[Lookup.scala 33:37]
  wire [4:0] _T_686 = _T_73 ? 5'h0 : _T_685; // @[Lookup.scala 33:37]
  wire [4:0] _T_687 = _T_71 ? 5'h0 : _T_686; // @[Lookup.scala 33:37]
  wire [4:0] _T_688 = _T_69 ? 5'h0 : _T_687; // @[Lookup.scala 33:37]
  wire [4:0] _T_689 = _T_67 ? 5'h0 : _T_688; // @[Lookup.scala 33:37]
  wire [4:0] _T_690 = _T_65 ? 5'h0 : _T_689; // @[Lookup.scala 33:37]
  wire [4:0] _T_691 = _T_63 ? 5'h0 : _T_690; // @[Lookup.scala 33:37]
  wire [4:0] _T_692 = _T_61 ? 5'h0 : _T_691; // @[Lookup.scala 33:37]
  wire [4:0] _T_693 = _T_59 ? 5'h0 : _T_692; // @[Lookup.scala 33:37]
  wire [4:0] _T_694 = _T_57 ? 5'h0 : _T_693; // @[Lookup.scala 33:37]
  wire [4:0] _T_695 = _T_55 ? 5'h0 : _T_694; // @[Lookup.scala 33:37]
  wire [4:0] _T_696 = _T_53 ? 5'h0 : _T_695; // @[Lookup.scala 33:37]
  wire [4:0] _T_697 = _T_51 ? 5'h0 : _T_696; // @[Lookup.scala 33:37]
  wire [4:0] _T_698 = _T_49 ? 5'h0 : _T_697; // @[Lookup.scala 33:37]
  wire [4:0] _T_699 = _T_47 ? 5'h0 : _T_698; // @[Lookup.scala 33:37]
  wire [4:0] _T_700 = _T_45 ? 5'h0 : _T_699; // @[Lookup.scala 33:37]
  wire [4:0] _T_701 = _T_43 ? 5'h0 : _T_700; // @[Lookup.scala 33:37]
  wire [4:0] _T_702 = _T_41 ? 5'h0 : _T_701; // @[Lookup.scala 33:37]
  wire [4:0] _T_703 = _T_39 ? 5'h0 : _T_702; // @[Lookup.scala 33:37]
  wire [4:0] _T_704 = _T_37 ? 5'h0 : _T_703; // @[Lookup.scala 33:37]
  wire [4:0] _T_705 = _T_35 ? 5'h0 : _T_704; // @[Lookup.scala 33:37]
  wire [4:0] _T_706 = _T_33 ? 5'h0 : _T_705; // @[Lookup.scala 33:37]
  wire [4:0] _T_707 = _T_31 ? 5'h0 : _T_706; // @[Lookup.scala 33:37]
  wire [4:0] _T_708 = _T_29 ? 5'h0 : _T_707; // @[Lookup.scala 33:37]
  wire [4:0] _T_709 = _T_27 ? 5'h0 : _T_708; // @[Lookup.scala 33:37]
  wire [4:0] _T_710 = _T_25 ? 5'h0 : _T_709; // @[Lookup.scala 33:37]
  wire [4:0] _T_711 = _T_23 ? 5'h0 : _T_710; // @[Lookup.scala 33:37]
  wire [4:0] lsuOp = _T_21 ? 5'h0 : _T_711; // @[Lookup.scala 33:37]
  wire [2:0] _T_737 = _T_109 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_738 = _T_107 ? 3'h4 : _T_737; // @[Lookup.scala 33:37]
  wire [2:0] _T_739 = _T_105 ? 3'h3 : _T_738; // @[Lookup.scala 33:37]
  wire [2:0] _T_740 = _T_103 ? 3'h5 : _T_739; // @[Lookup.scala 33:37]
  wire [2:0] _T_741 = _T_101 ? 3'h4 : _T_740; // @[Lookup.scala 33:37]
  wire [2:0] _T_742 = _T_99 ? 3'h3 : _T_741; // @[Lookup.scala 33:37]
  wire [2:0] _T_743 = _T_97 ? 3'h0 : _T_742; // @[Lookup.scala 33:37]
  wire [2:0] _T_744 = _T_95 ? 3'h0 : _T_743; // @[Lookup.scala 33:37]
  wire [2:0] _T_745 = _T_93 ? 3'h0 : _T_744; // @[Lookup.scala 33:37]
  wire [2:0] _T_746 = _T_91 ? 3'h0 : _T_745; // @[Lookup.scala 33:37]
  wire [2:0] _T_747 = _T_89 ? 3'h0 : _T_746; // @[Lookup.scala 33:37]
  wire [2:0] _T_748 = _T_87 ? 3'h0 : _T_747; // @[Lookup.scala 33:37]
  wire [2:0] _T_749 = _T_85 ? 3'h0 : _T_748; // @[Lookup.scala 33:37]
  wire [2:0] _T_750 = _T_83 ? 3'h0 : _T_749; // @[Lookup.scala 33:37]
  wire [2:0] _T_751 = _T_81 ? 3'h0 : _T_750; // @[Lookup.scala 33:37]
  wire [2:0] _T_752 = _T_79 ? 3'h0 : _T_751; // @[Lookup.scala 33:37]
  wire [2:0] _T_753 = _T_77 ? 3'h0 : _T_752; // @[Lookup.scala 33:37]
  wire [2:0] _T_754 = _T_75 ? 3'h0 : _T_753; // @[Lookup.scala 33:37]
  wire [2:0] _T_755 = _T_73 ? 3'h0 : _T_754; // @[Lookup.scala 33:37]
  wire [2:0] _T_756 = _T_71 ? 3'h0 : _T_755; // @[Lookup.scala 33:37]
  wire [2:0] _T_757 = _T_69 ? 3'h0 : _T_756; // @[Lookup.scala 33:37]
  wire [2:0] _T_758 = _T_67 ? 3'h0 : _T_757; // @[Lookup.scala 33:37]
  wire [2:0] _T_759 = _T_65 ? 3'h0 : _T_758; // @[Lookup.scala 33:37]
  wire [2:0] _T_760 = _T_63 ? 3'h0 : _T_759; // @[Lookup.scala 33:37]
  wire [2:0] _T_761 = _T_61 ? 3'h0 : _T_760; // @[Lookup.scala 33:37]
  wire [2:0] _T_762 = _T_59 ? 3'h0 : _T_761; // @[Lookup.scala 33:37]
  wire [2:0] _T_763 = _T_57 ? 3'h0 : _T_762; // @[Lookup.scala 33:37]
  wire [2:0] _T_764 = _T_55 ? 3'h0 : _T_763; // @[Lookup.scala 33:37]
  wire [2:0] _T_765 = _T_53 ? 3'h0 : _T_764; // @[Lookup.scala 33:37]
  wire [2:0] _T_766 = _T_51 ? 3'h0 : _T_765; // @[Lookup.scala 33:37]
  wire [2:0] _T_767 = _T_49 ? 3'h0 : _T_766; // @[Lookup.scala 33:37]
  wire [2:0] _T_768 = _T_47 ? 3'h0 : _T_767; // @[Lookup.scala 33:37]
  wire [2:0] _T_769 = _T_45 ? 3'h0 : _T_768; // @[Lookup.scala 33:37]
  wire [2:0] _T_770 = _T_43 ? 3'h0 : _T_769; // @[Lookup.scala 33:37]
  wire [2:0] _T_771 = _T_41 ? 3'h0 : _T_770; // @[Lookup.scala 33:37]
  wire [2:0] _T_772 = _T_39 ? 3'h0 : _T_771; // @[Lookup.scala 33:37]
  wire [2:0] _T_773 = _T_37 ? 3'h0 : _T_772; // @[Lookup.scala 33:37]
  wire [2:0] _T_774 = _T_35 ? 3'h0 : _T_773; // @[Lookup.scala 33:37]
  wire [2:0] _T_775 = _T_33 ? 3'h0 : _T_774; // @[Lookup.scala 33:37]
  wire [2:0] _T_776 = _T_31 ? 3'h0 : _T_775; // @[Lookup.scala 33:37]
  wire [2:0] _T_777 = _T_29 ? 3'h0 : _T_776; // @[Lookup.scala 33:37]
  wire [2:0] _T_778 = _T_27 ? 3'h0 : _T_777; // @[Lookup.scala 33:37]
  wire [2:0] _T_779 = _T_25 ? 3'h0 : _T_778; // @[Lookup.scala 33:37]
  wire [2:0] _T_780 = _T_23 ? 3'h0 : _T_779; // @[Lookup.scala 33:37]
  wire [2:0] csrOp = _T_21 ? 3'h0 : _T_780; // @[Lookup.scala 33:37]
  wire [3:0] _T_798 = _T_125 ? 4'h8 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_799 = _T_123 ? 4'h7 : _T_798; // @[Lookup.scala 33:37]
  wire [3:0] _T_800 = _T_121 ? 4'h6 : _T_799; // @[Lookup.scala 33:37]
  wire [3:0] _T_801 = _T_119 ? 4'h5 : _T_800; // @[Lookup.scala 33:37]
  wire [3:0] _T_802 = _T_117 ? 4'h4 : _T_801; // @[Lookup.scala 33:37]
  wire [3:0] _T_803 = _T_115 ? 4'h3 : _T_802; // @[Lookup.scala 33:37]
  wire [3:0] _T_804 = _T_113 ? 4'h2 : _T_803; // @[Lookup.scala 33:37]
  wire [3:0] _T_805 = _T_111 ? 4'h1 : _T_804; // @[Lookup.scala 33:37]
  wire [3:0] _T_806 = _T_109 ? 4'h0 : _T_805; // @[Lookup.scala 33:37]
  wire [3:0] _T_807 = _T_107 ? 4'h0 : _T_806; // @[Lookup.scala 33:37]
  wire [3:0] _T_808 = _T_105 ? 4'h0 : _T_807; // @[Lookup.scala 33:37]
  wire [3:0] _T_809 = _T_103 ? 4'h0 : _T_808; // @[Lookup.scala 33:37]
  wire [3:0] _T_810 = _T_101 ? 4'h0 : _T_809; // @[Lookup.scala 33:37]
  wire [3:0] _T_811 = _T_99 ? 4'h0 : _T_810; // @[Lookup.scala 33:37]
  wire [3:0] _T_812 = _T_97 ? 4'h0 : _T_811; // @[Lookup.scala 33:37]
  wire [3:0] _T_813 = _T_95 ? 4'h0 : _T_812; // @[Lookup.scala 33:37]
  wire [3:0] _T_814 = _T_93 ? 4'h0 : _T_813; // @[Lookup.scala 33:37]
  wire [3:0] _T_815 = _T_91 ? 4'h0 : _T_814; // @[Lookup.scala 33:37]
  wire [3:0] _T_816 = _T_89 ? 4'h0 : _T_815; // @[Lookup.scala 33:37]
  wire [3:0] _T_817 = _T_87 ? 4'h0 : _T_816; // @[Lookup.scala 33:37]
  wire [3:0] _T_818 = _T_85 ? 4'h0 : _T_817; // @[Lookup.scala 33:37]
  wire [3:0] _T_819 = _T_83 ? 4'h0 : _T_818; // @[Lookup.scala 33:37]
  wire [3:0] _T_820 = _T_81 ? 4'h0 : _T_819; // @[Lookup.scala 33:37]
  wire [3:0] _T_821 = _T_79 ? 4'h0 : _T_820; // @[Lookup.scala 33:37]
  wire [3:0] _T_822 = _T_77 ? 4'h0 : _T_821; // @[Lookup.scala 33:37]
  wire [3:0] _T_823 = _T_75 ? 4'h0 : _T_822; // @[Lookup.scala 33:37]
  wire [3:0] _T_824 = _T_73 ? 4'h0 : _T_823; // @[Lookup.scala 33:37]
  wire [3:0] _T_825 = _T_71 ? 4'h0 : _T_824; // @[Lookup.scala 33:37]
  wire [3:0] _T_826 = _T_69 ? 4'h0 : _T_825; // @[Lookup.scala 33:37]
  wire [3:0] _T_827 = _T_67 ? 4'h0 : _T_826; // @[Lookup.scala 33:37]
  wire [3:0] _T_828 = _T_65 ? 4'h0 : _T_827; // @[Lookup.scala 33:37]
  wire [3:0] _T_829 = _T_63 ? 4'h0 : _T_828; // @[Lookup.scala 33:37]
  wire [3:0] _T_830 = _T_61 ? 4'h0 : _T_829; // @[Lookup.scala 33:37]
  wire [3:0] _T_831 = _T_59 ? 4'h0 : _T_830; // @[Lookup.scala 33:37]
  wire [3:0] _T_832 = _T_57 ? 4'h0 : _T_831; // @[Lookup.scala 33:37]
  wire [3:0] _T_833 = _T_55 ? 4'h0 : _T_832; // @[Lookup.scala 33:37]
  wire [3:0] _T_834 = _T_53 ? 4'h0 : _T_833; // @[Lookup.scala 33:37]
  wire [3:0] _T_835 = _T_51 ? 4'h0 : _T_834; // @[Lookup.scala 33:37]
  wire [3:0] _T_836 = _T_49 ? 4'h0 : _T_835; // @[Lookup.scala 33:37]
  wire [3:0] _T_837 = _T_47 ? 4'h0 : _T_836; // @[Lookup.scala 33:37]
  wire [3:0] _T_838 = _T_45 ? 4'h0 : _T_837; // @[Lookup.scala 33:37]
  wire [3:0] _T_839 = _T_43 ? 4'h0 : _T_838; // @[Lookup.scala 33:37]
  wire [3:0] _T_840 = _T_41 ? 4'h0 : _T_839; // @[Lookup.scala 33:37]
  wire [3:0] _T_841 = _T_39 ? 4'h0 : _T_840; // @[Lookup.scala 33:37]
  wire [3:0] _T_842 = _T_37 ? 4'h0 : _T_841; // @[Lookup.scala 33:37]
  wire [3:0] _T_843 = _T_35 ? 4'h0 : _T_842; // @[Lookup.scala 33:37]
  wire [3:0] _T_844 = _T_33 ? 4'h0 : _T_843; // @[Lookup.scala 33:37]
  wire [3:0] _T_845 = _T_31 ? 4'h0 : _T_844; // @[Lookup.scala 33:37]
  wire [3:0] _T_846 = _T_29 ? 4'h0 : _T_845; // @[Lookup.scala 33:37]
  wire [3:0] _T_847 = _T_27 ? 4'h0 : _T_846; // @[Lookup.scala 33:37]
  wire [3:0] _T_848 = _T_25 ? 4'h0 : _T_847; // @[Lookup.scala 33:37]
  wire [3:0] _T_849 = _T_23 ? 4'h0 : _T_848; // @[Lookup.scala 33:37]
  wire [3:0] mduOp = _T_21 ? 4'h0 : _T_849; // @[Lookup.scala 33:37]
  wire [3:0] _T_850 = _T_159 ? 4'ha : 4'h5; // @[Lookup.scala 33:37]
  wire [3:0] _T_851 = _T_157 ? 4'h0 : _T_850; // @[Lookup.scala 33:37]
  wire [3:0] _T_852 = _T_155 ? 4'h4 : _T_851; // @[Lookup.scala 33:37]
  wire [3:0] _T_853 = _T_153 ? 4'h3 : _T_852; // @[Lookup.scala 33:37]
  wire [3:0] _T_854 = _T_151 ? 4'h2 : _T_853; // @[Lookup.scala 33:37]
  wire [3:0] _T_855 = _T_149 ? 4'h1 : _T_854; // @[Lookup.scala 33:37]
  wire [3:0] _T_856 = _T_147 ? 4'h9 : _T_855; // @[Lookup.scala 33:37]
  wire [3:0] _T_857 = _T_145 ? 4'h9 : _T_856; // @[Lookup.scala 33:37]
  wire [3:0] _T_858 = _T_143 ? 4'h9 : _T_857; // @[Lookup.scala 33:37]
  wire [3:0] _T_859 = _T_141 ? 4'h9 : _T_858; // @[Lookup.scala 33:37]
  wire [3:0] _T_860 = _T_139 ? 4'h9 : _T_859; // @[Lookup.scala 33:37]
  wire [3:0] _T_861 = _T_137 ? 4'h9 : _T_860; // @[Lookup.scala 33:37]
  wire [3:0] _T_862 = _T_135 ? 4'h9 : _T_861; // @[Lookup.scala 33:37]
  wire [3:0] _T_863 = _T_133 ? 4'h9 : _T_862; // @[Lookup.scala 33:37]
  wire [3:0] _T_864 = _T_131 ? 4'h9 : _T_863; // @[Lookup.scala 33:37]
  wire [3:0] _T_865 = _T_129 ? 4'h9 : _T_864; // @[Lookup.scala 33:37]
  wire [3:0] _T_866 = _T_127 ? 4'h9 : _T_865; // @[Lookup.scala 33:37]
  wire [3:0] _T_867 = _T_125 ? 4'h0 : _T_866; // @[Lookup.scala 33:37]
  wire [3:0] _T_868 = _T_123 ? 4'h0 : _T_867; // @[Lookup.scala 33:37]
  wire [3:0] _T_869 = _T_121 ? 4'h0 : _T_868; // @[Lookup.scala 33:37]
  wire [3:0] _T_870 = _T_119 ? 4'h0 : _T_869; // @[Lookup.scala 33:37]
  wire [3:0] _T_871 = _T_117 ? 4'h0 : _T_870; // @[Lookup.scala 33:37]
  wire [3:0] _T_872 = _T_115 ? 4'h0 : _T_871; // @[Lookup.scala 33:37]
  wire [3:0] _T_873 = _T_113 ? 4'h0 : _T_872; // @[Lookup.scala 33:37]
  wire [3:0] _T_874 = _T_111 ? 4'h0 : _T_873; // @[Lookup.scala 33:37]
  wire [3:0] _T_875 = _T_109 ? 4'h0 : _T_874; // @[Lookup.scala 33:37]
  wire [3:0] _T_876 = _T_107 ? 4'h0 : _T_875; // @[Lookup.scala 33:37]
  wire [3:0] _T_877 = _T_105 ? 4'h0 : _T_876; // @[Lookup.scala 33:37]
  wire [3:0] _T_878 = _T_103 ? 4'h0 : _T_877; // @[Lookup.scala 33:37]
  wire [3:0] _T_879 = _T_101 ? 4'h0 : _T_878; // @[Lookup.scala 33:37]
  wire [3:0] _T_880 = _T_99 ? 4'h0 : _T_879; // @[Lookup.scala 33:37]
  wire [3:0] _T_881 = _T_97 ? 4'h0 : _T_880; // @[Lookup.scala 33:37]
  wire [3:0] _T_882 = _T_95 ? 4'h0 : _T_881; // @[Lookup.scala 33:37]
  wire [3:0] _T_883 = _T_93 ? 4'h9 : _T_882; // @[Lookup.scala 33:37]
  wire [3:0] _T_884 = _T_91 ? 4'h9 : _T_883; // @[Lookup.scala 33:37]
  wire [3:0] _T_885 = _T_89 ? 4'h9 : _T_884; // @[Lookup.scala 33:37]
  wire [3:0] _T_886 = _T_87 ? 4'h8 : _T_885; // @[Lookup.scala 33:37]
  wire [3:0] _T_887 = _T_85 ? 4'h8 : _T_886; // @[Lookup.scala 33:37]
  wire [3:0] _T_888 = _T_83 ? 4'h8 : _T_887; // @[Lookup.scala 33:37]
  wire [3:0] _T_889 = _T_81 ? 4'h8 : _T_888; // @[Lookup.scala 33:37]
  wire [3:0] _T_890 = _T_79 ? 4'h8 : _T_889; // @[Lookup.scala 33:37]
  wire [3:0] _T_891 = _T_77 ? 4'h0 : _T_890; // @[Lookup.scala 33:37]
  wire [3:0] _T_892 = _T_75 ? 4'h0 : _T_891; // @[Lookup.scala 33:37]
  wire [3:0] _T_893 = _T_73 ? 4'h0 : _T_892; // @[Lookup.scala 33:37]
  wire [3:0] _T_894 = _T_71 ? 4'h0 : _T_893; // @[Lookup.scala 33:37]
  wire [3:0] _T_895 = _T_69 ? 4'h0 : _T_894; // @[Lookup.scala 33:37]
  wire [3:0] _T_896 = _T_67 ? 4'h0 : _T_895; // @[Lookup.scala 33:37]
  wire [3:0] _T_897 = _T_65 ? 4'h0 : _T_896; // @[Lookup.scala 33:37]
  wire [3:0] _T_898 = _T_63 ? 4'h0 : _T_897; // @[Lookup.scala 33:37]
  wire [3:0] _T_899 = _T_61 ? 4'h0 : _T_898; // @[Lookup.scala 33:37]
  wire [3:0] _T_900 = _T_59 ? 4'h0 : _T_899; // @[Lookup.scala 33:37]
  wire [3:0] _T_901 = _T_57 ? 4'h0 : _T_900; // @[Lookup.scala 33:37]
  wire [3:0] _T_902 = _T_55 ? 4'h0 : _T_901; // @[Lookup.scala 33:37]
  wire [3:0] _T_903 = _T_53 ? 4'h0 : _T_902; // @[Lookup.scala 33:37]
  wire [3:0] _T_904 = _T_51 ? 4'h0 : _T_903; // @[Lookup.scala 33:37]
  wire [3:0] _T_905 = _T_49 ? 4'h0 : _T_904; // @[Lookup.scala 33:37]
  wire [3:0] _T_906 = _T_47 ? 4'h0 : _T_905; // @[Lookup.scala 33:37]
  wire [3:0] _T_907 = _T_45 ? 4'h0 : _T_906; // @[Lookup.scala 33:37]
  wire [3:0] _T_908 = _T_43 ? 4'h0 : _T_907; // @[Lookup.scala 33:37]
  wire [3:0] _T_909 = _T_41 ? 4'h0 : _T_908; // @[Lookup.scala 33:37]
  wire [3:0] _T_910 = _T_39 ? 4'h0 : _T_909; // @[Lookup.scala 33:37]
  wire [3:0] _T_911 = _T_37 ? 4'h0 : _T_910; // @[Lookup.scala 33:37]
  wire [3:0] _T_912 = _T_35 ? 4'h0 : _T_911; // @[Lookup.scala 33:37]
  wire [3:0] _T_913 = _T_33 ? 4'h0 : _T_912; // @[Lookup.scala 33:37]
  wire [3:0] _T_914 = _T_31 ? 4'h0 : _T_913; // @[Lookup.scala 33:37]
  wire [3:0] _T_915 = _T_29 ? 4'h0 : _T_914; // @[Lookup.scala 33:37]
  wire [3:0] _T_916 = _T_27 ? 4'h0 : _T_915; // @[Lookup.scala 33:37]
  wire [3:0] _T_917 = _T_25 ? 4'h0 : _T_916; // @[Lookup.scala 33:37]
  wire [3:0] _T_918 = _T_23 ? 4'h0 : _T_917; // @[Lookup.scala 33:37]
  wire [3:0] excType = _T_21 ? 4'h0 : _T_918; // @[Lookup.scala 33:37]
  wire  isJump = branchFlag == 3'h1; // @[Decoder.scala 74:32]
  wire [20:0] _T_920 = {inst[31],inst[19:12],inst[20],inst[30:21],1'h0}; // @[Decoder.scala 75:48]
  wire [31:0] _GEN_1 = {{11{_T_920[20]}},_T_920}; // @[Decoder.scala 75:41]
  wire [31:0] targetJAL = $signed(io_fetch_pc) + $signed(_GEN_1); // @[Decoder.scala 75:56]
  wire [11:0] _T_925 = inst[31:20]; // @[Decoder.scala 76:49]
  wire [31:0] _GEN_2 = {{20{_T_925[11]}},_T_925}; // @[Decoder.scala 76:42]
  wire [31:0] sumR1immI = $signed(io_read1_data) + $signed(_GEN_2); // @[Decoder.scala 76:42]
  wire [31:0] targetJALR = {sumR1immI[31:1],1'h0}; // @[Cat.scala 30:58]
  wire [31:0] targetJ = regEn1 ? targetJALR : targetJAL; // @[Decoder.scala 78:24]
  wire [12:0] _T_930 = {inst[31],inst[7],inst[30:25],inst[11:8],1'h0}; // @[Decoder.scala 79:48]
  wire [31:0] _GEN_3 = {{19{_T_930[12]}},_T_930}; // @[Decoder.scala 79:41]
  wire [31:0] targetB = $signed(io_fetch_pc) + $signed(_GEN_3); // @[Decoder.scala 79:56]
  wire  _T_934 = io_read1_data == io_read2_data; // @[Decoder.scala 83:31]
  wire  _T_935 = io_read1_data != io_read2_data; // @[Decoder.scala 84:31]
  wire  _T_938 = $signed(io_read1_data) < $signed(io_read2_data); // @[Decoder.scala 85:38]
  wire  _T_941 = $signed(io_read1_data) >= $signed(io_read2_data); // @[Decoder.scala 86:38]
  wire  _T_942 = io_read1_data < io_read2_data; // @[Decoder.scala 87:31]
  wire  _T_943 = io_read1_data >= io_read2_data; // @[Decoder.scala 88:31]
  wire  _T_944 = 3'h7 == branchFlag; // @[Mux.scala 68:19]
  wire  _T_945 = _T_944 & _T_943; // @[Mux.scala 68:16]
  wire  _T_946 = 3'h6 == branchFlag; // @[Mux.scala 68:19]
  wire  _T_947 = _T_946 ? _T_942 : _T_945; // @[Mux.scala 68:16]
  wire  _T_948 = 3'h5 == branchFlag; // @[Mux.scala 68:19]
  wire  _T_949 = _T_948 ? _T_941 : _T_947; // @[Mux.scala 68:16]
  wire  _T_950 = 3'h4 == branchFlag; // @[Mux.scala 68:19]
  wire  _T_951 = _T_950 ? _T_938 : _T_949; // @[Mux.scala 68:16]
  wire  _T_952 = 3'h3 == branchFlag; // @[Mux.scala 68:19]
  wire  _T_953 = _T_952 ? _T_935 : _T_951; // @[Mux.scala 68:16]
  wire  _T_954 = 3'h2 == branchFlag; // @[Mux.scala 68:19]
  wire  _T_955 = _T_954 ? _T_934 : _T_953; // @[Mux.scala 68:16]
  wire  _T_956 = 3'h1 == branchFlag; // @[Mux.scala 68:19]
  wire  branchTaken = _T_956 | _T_955; // @[Mux.scala 68:16]
  wire  _T_957 = branchFlag == 3'h0; // @[Decoder.scala 90:38]
  wire [31:0] _T_958 = isJump ? targetJ : targetB; // @[Decoder.scala 91:26]
  wire [31:0] branchTarget = _T_957 ? 32'h0 : _T_958; // @[Decoder.scala 90:26]
  wire  _T_959 = io_fetch_taken != branchTaken; // @[Decoder.scala 92:36]
  wire  _T_960 = io_fetch_target != branchTarget; // @[Decoder.scala 93:53]
  wire  _T_961 = branchTaken & _T_960; // @[Decoder.scala 93:34]
  wire  branchMiss = _T_959 | _T_961; // @[Decoder.scala 92:52]
  wire [31:0] _T_963 = io_fetch_pc + 32'h4; // @[Decoder.scala 94:64]
  wire  _T_965 = branchTarget[1:0] != 2'h0; // @[Decoder.scala 96:59]
  wire  addrFault = branchTaken & _T_965; // @[Decoder.scala 95:33]
  wire  _T_966 = rd == 5'h0; // @[Decoder.scala 100:23]
  wire [2:0] _T_967 = _T_966 ? 3'h2 : 3'h3; // @[Decoder.scala 100:19]
  wire  _T_968 = rs1 == 5'h0; // @[Decoder.scala 101:24]
  wire [2:0] _T_969 = _T_968 ? 3'h1 : 3'h4; // @[Decoder.scala 101:19]
  wire [2:0] _T_971 = _T_968 ? 3'h1 : 3'h5; // @[Decoder.scala 102:19]
  wire  _T_972 = 3'h5 == csrOp; // @[Mux.scala 68:19]
  wire [2:0] _T_973 = _T_972 ? _T_971 : 3'h0; // @[Mux.scala 68:16]
  wire  _T_974 = 3'h4 == csrOp; // @[Mux.scala 68:19]
  wire [2:0] _T_975 = _T_974 ? _T_969 : _T_973; // @[Mux.scala 68:16]
  wire  _T_976 = 3'h3 == csrOp; // @[Mux.scala 68:19]
  wire [2:0] csrActOp = _T_976 ? _T_967 : _T_975; // @[Mux.scala 68:16]
  wire  _T_977 = csrActOp == 3'h0; // @[Decoder.scala 104:32]
  wire [31:0] _T_978 = regEn1 ? io_read1_data : {{27'd0}, rs1}; // @[Decoder.scala 105:22]
  wire [3:0] _T_979 = addrFault ? 4'h7 : excType; // @[Decoder.scala 109:24]
  wire [3:0] exceptType = io_fetch_pageFault ? 4'h6 : _T_979; // @[Decoder.scala 108:24]
  wire  _T_980 = exceptType == 4'h5; // @[Decoder.scala 114:34]
  wire  _T_981 = exceptType == 4'h6; // @[Decoder.scala 114:62]
  wire  illegalFetch = _T_980 | _T_981; // @[Decoder.scala 114:48]
  wire  _T_982 = ~io_stallId; // @[Decoder.scala 120:18]
  wire  _T_983 = ~addrFault; // @[Decoder.scala 120:33]
  wire  _T_984 = _T_982 & _T_983; // @[Decoder.scala 120:30]
  wire [11:0] _T_989 = {inst[31:25],rd}; // @[Decoder.scala 60:27]
  wire [31:0] _T_990 = {inst[31:12],12'h0}; // @[Decoder.scala 61:27]
  wire [5:0] _T_991 = {1'b0,$signed(rs2)}; // @[Decoder.scala 62:26]
  wire  _T_993 = 4'h8 == aluSrc1; // @[Mux.scala 68:19]
  wire [3:0] _T_994 = _T_993 ? $signed(4'sh4) : $signed(4'sh0); // @[Mux.scala 68:16]
  wire  _T_995 = 4'h7 == aluSrc1; // @[Mux.scala 68:19]
  wire [31:0] _T_996 = _T_995 ? $signed(io_fetch_pc) : $signed({{28{_T_994[3]}},_T_994}); // @[Mux.scala 68:16]
  wire  _T_997 = 4'h6 == aluSrc1; // @[Mux.scala 68:19]
  wire [31:0] _T_998 = _T_997 ? $signed({{26{_T_991[5]}},_T_991}) : $signed(_T_996); // @[Mux.scala 68:16]
  wire  _T_999 = 4'h5 == aluSrc1; // @[Mux.scala 68:19]
  wire [31:0] _T_1000 = _T_999 ? $signed(_T_990) : $signed(_T_998); // @[Mux.scala 68:16]
  wire  _T_1001 = 4'h4 == aluSrc1; // @[Mux.scala 68:19]
  wire [31:0] _T_1002 = _T_1001 ? $signed({{20{_T_989[11]}},_T_989}) : $signed(_T_1000); // @[Mux.scala 68:16]
  wire  _T_1003 = 4'h3 == aluSrc1; // @[Mux.scala 68:19]
  wire [31:0] _T_1004 = _T_1003 ? $signed({{20{_T_925[11]}},_T_925}) : $signed(_T_1002); // @[Mux.scala 68:16]
  wire  _T_1005 = 4'h2 == aluSrc1; // @[Mux.scala 68:19]
  wire [31:0] _T_1006 = _T_1005 ? $signed(io_read2_data) : $signed(_T_1004); // @[Mux.scala 68:16]
  wire  _T_1007 = 4'h1 == aluSrc1; // @[Mux.scala 68:19]
  wire  _T_1017 = 4'h8 == aluSrc2; // @[Mux.scala 68:19]
  wire [3:0] _T_1018 = _T_1017 ? $signed(4'sh4) : $signed(4'sh0); // @[Mux.scala 68:16]
  wire  _T_1019 = 4'h7 == aluSrc2; // @[Mux.scala 68:19]
  wire [31:0] _T_1020 = _T_1019 ? $signed(io_fetch_pc) : $signed({{28{_T_1018[3]}},_T_1018}); // @[Mux.scala 68:16]
  wire  _T_1021 = 4'h6 == aluSrc2; // @[Mux.scala 68:19]
  wire [31:0] _T_1022 = _T_1021 ? $signed({{26{_T_991[5]}},_T_991}) : $signed(_T_1020); // @[Mux.scala 68:16]
  wire  _T_1023 = 4'h5 == aluSrc2; // @[Mux.scala 68:19]
  wire [31:0] _T_1024 = _T_1023 ? $signed(_T_990) : $signed(_T_1022); // @[Mux.scala 68:16]
  wire  _T_1025 = 4'h4 == aluSrc2; // @[Mux.scala 68:19]
  wire [31:0] _T_1026 = _T_1025 ? $signed({{20{_T_989[11]}},_T_989}) : $signed(_T_1024); // @[Mux.scala 68:16]
  wire  _T_1027 = 4'h3 == aluSrc2; // @[Mux.scala 68:19]
  wire [31:0] _T_1028 = _T_1027 ? $signed({{20{_T_925[11]}},_T_925}) : $signed(_T_1026); // @[Mux.scala 68:16]
  wire  _T_1029 = 4'h2 == aluSrc2; // @[Mux.scala 68:19]
  wire [31:0] _T_1030 = _T_1029 ? $signed(io_read2_data) : $signed(_T_1028); // @[Mux.scala 68:16]
  wire  _T_1031 = 4'h1 == aluSrc2; // @[Mux.scala 68:19]
  assign io_flushIf = _T_984 & branchMiss; // @[Decoder.scala 120:15]
  assign io_flushPc = branchTaken ? branchTarget : _T_963; // @[Decoder.scala 121:15]
  assign io_read1_en = _T_21 | _T_228; // @[Decoder.scala 124:17]
  assign io_read1_addr = inst[19:15]; // @[Decoder.scala 125:17]
  assign io_read2_en = _T_21 | _T_297; // @[Decoder.scala 126:17]
  assign io_read2_addr = inst[24:20]; // @[Decoder.scala 127:17]
  assign io_branch_branch = branchFlag != 3'h0; // @[Decoder.scala 130:21]
  assign io_branch_jump = branchFlag == 3'h1; // @[Decoder.scala 131:21]
  assign io_branch_taken = _T_956 | _T_955; // @[Decoder.scala 132:21]
  assign io_branch_index = io_fetch_predIndex; // @[Decoder.scala 133:21]
  assign io_branch_pc = io_fetch_pc; // @[Decoder.scala 134:21]
  assign io_branch_target = _T_957 ? 32'h0 : _T_958; // @[Decoder.scala 135:21]
  assign io_decoder_aluOp = _T_21 ? 4'h0 : _T_573; // @[Decoder.scala 139:25]
  assign io_decoder_opr1 = _T_1007 ? $signed(io_read1_data) : $signed(_T_1006); // @[Decoder.scala 140:25]
  assign io_decoder_opr2 = _T_1031 ? $signed(io_read1_data) : $signed(_T_1030); // @[Decoder.scala 141:25]
  assign io_decoder_mduOp = illegalFetch ? 4'h0 : mduOp; // @[Decoder.scala 142:25]
  assign io_decoder_lsuOp = illegalFetch ? 5'h0 : lsuOp; // @[Decoder.scala 144:25]
  assign io_decoder_lsuData = io_read2_data; // @[Decoder.scala 145:25]
  assign io_decoder_regWen = _T_21 | _T_366; // @[Decoder.scala 147:25]
  assign io_decoder_regWaddr = inst[11:7]; // @[Decoder.scala 148:25]
  assign io_decoder_csrOp = illegalFetch ? 3'h0 : csrActOp; // @[Decoder.scala 150:25]
  assign io_decoder_csrAddr = inst[31:20]; // @[Decoder.scala 151:25]
  assign io_decoder_csrData = _T_977 ? 32'h0 : _T_978; // @[Decoder.scala 152:25]
  assign io_decoder_excType = io_fetch_pageFault ? 4'h6 : _T_979; // @[Decoder.scala 154:25]
  assign io_decoder_excValue = addrFault ? branchTarget : 32'h0; // @[Decoder.scala 155:25]
  assign io_decoder_valid = io_fetch_valid; // @[Decoder.scala 157:25]
  assign io_decoder_inst = _T ? 32'h13 : _T_1; // @[Decoder.scala 158:25]
  assign io_decoder_currentPc = io_fetch_pc; // @[Decoder.scala 159:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stallDelay = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  lastInst = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    stallDelay <= io_stallId;
    if (_T_2) begin
      lastInst <= io_inst;
    end
  end
endmodule
module MidStage_1(
  input         clock,
  input         reset,
  input         io_flush,
  input         io_stallPrev,
  input         io_stallNext,
  input  [3:0]  io_prev_aluOp,
  input  [31:0] io_prev_opr1,
  input  [31:0] io_prev_opr2,
  input  [3:0]  io_prev_mduOp,
  input  [4:0]  io_prev_lsuOp,
  input  [31:0] io_prev_lsuData,
  input         io_prev_regWen,
  input  [4:0]  io_prev_regWaddr,
  input  [2:0]  io_prev_csrOp,
  input  [11:0] io_prev_csrAddr,
  input  [31:0] io_prev_csrData,
  input  [3:0]  io_prev_excType,
  input  [31:0] io_prev_excValue,
  input         io_prev_valid,
  input  [31:0] io_prev_inst,
  input  [31:0] io_prev_currentPc,
  output [3:0]  io_next_aluOp,
  output [31:0] io_next_opr1,
  output [31:0] io_next_opr2,
  output [3:0]  io_next_mduOp,
  output [4:0]  io_next_lsuOp,
  output [31:0] io_next_lsuData,
  output        io_next_regWen,
  output [4:0]  io_next_regWaddr,
  output [2:0]  io_next_csrOp,
  output [11:0] io_next_csrAddr,
  output [31:0] io_next_csrData,
  output [3:0]  io_next_excType,
  output [31:0] io_next_excValue,
  output        io_next_valid,
  output [31:0] io_next_inst,
  output [31:0] io_next_currentPc
);
  reg [3:0] ff_aluOp; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_0;
  reg [31:0] ff_opr1; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_1;
  reg [31:0] ff_opr2; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_2;
  reg [3:0] ff_mduOp; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_3;
  reg [4:0] ff_lsuOp; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_4;
  reg [31:0] ff_lsuData; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_5;
  reg  ff_regWen; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_6;
  reg [4:0] ff_regWaddr; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_7;
  reg [2:0] ff_csrOp; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_8;
  reg [11:0] ff_csrAddr; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_9;
  reg [31:0] ff_csrData; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_10;
  reg [3:0] ff_excType; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_11;
  reg [31:0] ff_excValue; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_12;
  reg  ff_valid; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_13;
  reg [31:0] ff_inst; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_14;
  reg [31:0] ff_currentPc; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_15;
  wire  _T_1 = ~io_stallNext; // @[MidStage.scala 21:38]
  wire  _T_2 = io_stallPrev & _T_1; // @[MidStage.scala 21:35]
  wire  _T_3 = io_flush | _T_2; // @[MidStage.scala 21:18]
  wire  _T_5 = ~io_stallPrev; // @[MidStage.scala 23:15]
  assign io_next_aluOp = ff_aluOp; // @[MidStage.scala 27:11]
  assign io_next_opr1 = ff_opr1; // @[MidStage.scala 27:11]
  assign io_next_opr2 = ff_opr2; // @[MidStage.scala 27:11]
  assign io_next_mduOp = ff_mduOp; // @[MidStage.scala 27:11]
  assign io_next_lsuOp = ff_lsuOp; // @[MidStage.scala 27:11]
  assign io_next_lsuData = ff_lsuData; // @[MidStage.scala 27:11]
  assign io_next_regWen = ff_regWen; // @[MidStage.scala 27:11]
  assign io_next_regWaddr = ff_regWaddr; // @[MidStage.scala 27:11]
  assign io_next_csrOp = ff_csrOp; // @[MidStage.scala 27:11]
  assign io_next_csrAddr = ff_csrAddr; // @[MidStage.scala 27:11]
  assign io_next_csrData = ff_csrData; // @[MidStage.scala 27:11]
  assign io_next_excType = ff_excType; // @[MidStage.scala 27:11]
  assign io_next_excValue = ff_excValue; // @[MidStage.scala 27:11]
  assign io_next_valid = ff_valid; // @[MidStage.scala 27:11]
  assign io_next_inst = ff_inst; // @[MidStage.scala 27:11]
  assign io_next_currentPc = ff_currentPc; // @[MidStage.scala 27:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff_aluOp = _RAND_0[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ff_opr1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ff_opr2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ff_mduOp = _RAND_3[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ff_lsuOp = _RAND_4[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ff_lsuData = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ff_regWen = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ff_regWaddr = _RAND_7[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ff_csrOp = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  ff_csrAddr = _RAND_9[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  ff_csrData = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  ff_excType = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  ff_excValue = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  ff_valid = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  ff_inst = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  ff_currentPc = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ff_aluOp <= 4'h0;
    end else if (_T_3) begin
      ff_aluOp <= 4'h0;
    end else if (_T_5) begin
      ff_aluOp <= io_prev_aluOp;
    end
    if (reset) begin
      ff_opr1 <= 32'h0;
    end else if (_T_3) begin
      ff_opr1 <= 32'h0;
    end else if (_T_5) begin
      ff_opr1 <= io_prev_opr1;
    end
    if (reset) begin
      ff_opr2 <= 32'h0;
    end else if (_T_3) begin
      ff_opr2 <= 32'h0;
    end else if (_T_5) begin
      ff_opr2 <= io_prev_opr2;
    end
    if (reset) begin
      ff_mduOp <= 4'h0;
    end else if (_T_3) begin
      ff_mduOp <= 4'h0;
    end else if (_T_5) begin
      ff_mduOp <= io_prev_mduOp;
    end
    if (reset) begin
      ff_lsuOp <= 5'h0;
    end else if (_T_3) begin
      ff_lsuOp <= 5'h0;
    end else if (_T_5) begin
      ff_lsuOp <= io_prev_lsuOp;
    end
    if (reset) begin
      ff_lsuData <= 32'h0;
    end else if (_T_3) begin
      ff_lsuData <= 32'h0;
    end else if (_T_5) begin
      ff_lsuData <= io_prev_lsuData;
    end
    if (reset) begin
      ff_regWen <= 1'h0;
    end else if (_T_3) begin
      ff_regWen <= 1'h0;
    end else if (_T_5) begin
      ff_regWen <= io_prev_regWen;
    end
    if (reset) begin
      ff_regWaddr <= 5'h0;
    end else if (_T_3) begin
      ff_regWaddr <= 5'h0;
    end else if (_T_5) begin
      ff_regWaddr <= io_prev_regWaddr;
    end
    if (reset) begin
      ff_csrOp <= 3'h0;
    end else if (_T_3) begin
      ff_csrOp <= 3'h0;
    end else if (_T_5) begin
      ff_csrOp <= io_prev_csrOp;
    end
    if (reset) begin
      ff_csrAddr <= 12'h0;
    end else if (_T_3) begin
      ff_csrAddr <= 12'h0;
    end else if (_T_5) begin
      ff_csrAddr <= io_prev_csrAddr;
    end
    if (reset) begin
      ff_csrData <= 32'h0;
    end else if (_T_3) begin
      ff_csrData <= 32'h0;
    end else if (_T_5) begin
      ff_csrData <= io_prev_csrData;
    end
    if (reset) begin
      ff_excType <= 4'h0;
    end else if (_T_3) begin
      ff_excType <= 4'h0;
    end else if (_T_5) begin
      ff_excType <= io_prev_excType;
    end
    if (reset) begin
      ff_excValue <= 32'h0;
    end else if (_T_3) begin
      ff_excValue <= 32'h0;
    end else if (_T_5) begin
      ff_excValue <= io_prev_excValue;
    end
    if (reset) begin
      ff_valid <= 1'h0;
    end else if (_T_3) begin
      ff_valid <= 1'h0;
    end else if (_T_5) begin
      ff_valid <= io_prev_valid;
    end
    if (reset) begin
      ff_inst <= 32'h0;
    end else if (_T_3) begin
      ff_inst <= 32'h0;
    end else if (_T_5) begin
      ff_inst <= io_prev_inst;
    end
    if (reset) begin
      ff_currentPc <= 32'h0;
    end else if (_T_3) begin
      ff_currentPc <= 32'h0;
    end else if (_T_5) begin
      ff_currentPc <= io_prev_currentPc;
    end
  end
endmodule
module Multiplier(
  input         clock,
  input         reset,
  input         io_en,
  input         io_flush,
  output        io_done,
  input  [31:0] io_opr1,
  input  [31:0] io_opr2,
  output [63:0] io_result
);
  wire [63:0] result = io_opr1 * io_opr2; // @[Multiplier.scala 23:25]
  reg  en; // @[Multiplier.scala 30:26]
  reg [31:0] _RAND_0;
  reg [63:0] data; // @[Reg.scala 15:16]
  reg [63:0] _RAND_1;
  assign io_done = en; // @[Multiplier.scala 38:18]
  assign io_result = data; // @[Multiplier.scala 39:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  en = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {2{`RANDOM}};
  data = _RAND_1[63:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      en <= 1'h0;
    end else if (io_flush) begin
      en <= 1'h0;
    end else begin
      en <= io_en;
    end
    if (io_en) begin
      data <= result;
    end
  end
endmodule
module Divider(
  input         clock,
  input         reset,
  input         io_en,
  input         io_flush,
  output        io_divZero,
  output        io_done,
  input  [31:0] io_divident,
  input  [31:0] io_divisor,
  output [31:0] io_quotient,
  output [31:0] io_remainder
);
  reg [1:0] state; // @[Divider.scala 27:22]
  reg [31:0] _RAND_0;
  reg [64:0] result; // @[Divider.scala 31:30]
  reg [95:0] _RAND_1;
  reg [3:0] counter; // @[Divider.scala 33:30]
  reg [31:0] _RAND_2;
  reg  isDiv0; // @[Divider.scala 35:30]
  reg [31:0] _RAND_3;
  reg [31:0] lastDivident; // @[Divider.scala 37:30]
  reg [31:0] _RAND_4;
  reg [31:0] lastDivisor; // @[Divider.scala 38:30]
  reg [31:0] _RAND_5;
  reg [64:0] divisor; // @[Divider.scala 41:28]
  reg [95:0] _RAND_6;
  wire [63:0] minDivisor = divisor[64:1]; // @[Divider.scala 43:29]
  wire [64:0] _GEN_41 = {{1'd0}, minDivisor}; // @[Divider.scala 45:29]
  wire [64:0] maxDivisor = divisor + _GEN_41; // @[Divider.scala 45:29]
  wire  _T_1 = lastDivident != io_divident; // @[Divider.scala 47:34]
  wire  _T_2 = lastDivisor != io_divisor; // @[Divider.scala 48:33]
  wire  startFlag = _T_1 | _T_2; // @[Divider.scala 47:50]
  wire  _T_3 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = io_divisor == 32'h0; // @[Divider.scala 64:30]
  wire [64:0] _T_6 = {32'h0,io_divident,1'h0}; // @[Cat.scala 30:58]
  wire [64:0] _T_8 = {1'h0,io_divisor,32'h0}; // @[Cat.scala 30:58]
  wire [64:0] _GEN_2 = _T_4 ? result : _T_6; // @[Divider.scala 64:39]
  wire [64:0] _GEN_9 = startFlag ? _GEN_2 : result; // @[Divider.scala 59:28]
  wire [64:0] _GEN_16 = io_en ? _GEN_9 : result; // @[Divider.scala 58:22]
  wire  _T_9 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = result >= maxDivisor; // @[Divider.scala 82:22]
  wire [64:0] _T_12 = result - maxDivisor; // @[Divider.scala 83:30]
  wire [66:0] _T_13 = {_T_12, 2'h0}; // @[Divider.scala 83:44]
  wire [66:0] _T_14 = _T_13 | 67'h3; // @[Divider.scala 83:50]
  wire  _T_15 = result < maxDivisor; // @[Divider.scala 84:29]
  wire  _T_16 = result >= divisor; // @[Divider.scala 84:52]
  wire  _T_17 = _T_15 & _T_16; // @[Divider.scala 84:42]
  wire [64:0] _T_19 = result - divisor; // @[Divider.scala 85:30]
  wire [66:0] _T_20 = {_T_19, 2'h0}; // @[Divider.scala 85:41]
  wire [66:0] _T_21 = _T_20 | 67'h2; // @[Divider.scala 85:47]
  wire  _T_22 = result < divisor; // @[Divider.scala 86:29]
  wire  _T_23 = result >= _GEN_41; // @[Divider.scala 86:49]
  wire  _T_24 = _T_22 & _T_23; // @[Divider.scala 86:39]
  wire [64:0] _T_26 = result - _GEN_41; // @[Divider.scala 87:30]
  wire [66:0] _T_27 = {_T_26, 2'h0}; // @[Divider.scala 87:44]
  wire [66:0] _T_28 = _T_27 | 67'h1; // @[Divider.scala 87:50]
  wire [66:0] _T_29 = {result, 2'h0}; // @[Divider.scala 89:28]
  wire [66:0] _GEN_19 = _T_24 ? _T_28 : _T_29; // @[Divider.scala 86:64]
  wire [66:0] _GEN_20 = _T_17 ? _T_21 : _GEN_19; // @[Divider.scala 84:64]
  wire [66:0] _GEN_21 = _T_10 ? _T_14 : _GEN_20; // @[Divider.scala 82:37]
  wire [3:0] _T_31 = counter + 4'h1; // @[Divider.scala 92:28]
  wire  _T_32 = counter == 4'hf; // @[Divider.scala 93:23]
  wire  _T_33 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [66:0] _GEN_24 = _T_9 ? _GEN_21 : {{2'd0}, result}; // @[Conditional.scala 39:67]
  wire [66:0] _GEN_31 = _T_3 ? {{2'd0}, _GEN_16} : _GEN_24; // @[Conditional.scala 40:58]
  wire [66:0] _GEN_35 = io_flush ? 67'h0 : _GEN_31; // @[Divider.scala 51:19]
  assign io_divZero = isDiv0; // @[Divider.scala 102:17]
  assign io_done = state == 2'h2; // @[Divider.scala 103:17]
  assign io_quotient = result[31:0]; // @[Divider.scala 104:17]
  assign io_remainder = result[64:33]; // @[Divider.scala 105:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {3{`RANDOM}};
  result = _RAND_1[64:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  counter = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  isDiv0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  lastDivident = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  lastDivisor = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {3{`RANDOM}};
  divisor = _RAND_6[64:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (io_flush) begin
      state <= 2'h0;
    end else if (_T_3) begin
      if (io_en) begin
        if (startFlag) begin
          if (_T_4) begin
            state <= 2'h2;
          end else begin
            state <= 2'h1;
          end
        end else begin
          state <= 2'h2;
        end
      end
    end else if (_T_9) begin
      if (_T_32) begin
        state <= 2'h2;
      end
    end else if (_T_33) begin
      state <= 2'h0;
    end
    if (reset) begin
      result <= 65'h0;
    end else begin
      result <= _GEN_35[64:0];
    end
    if (reset) begin
      counter <= 4'h0;
    end else if (!(io_flush)) begin
      if (_T_3) begin
        if (io_en) begin
          if (startFlag) begin
            if (!(_T_4)) begin
              counter <= 4'h0;
            end
          end
        end
      end else if (_T_9) begin
        counter <= _T_31;
      end
    end
    if (reset) begin
      isDiv0 <= 1'h0;
    end else if (io_flush) begin
      isDiv0 <= 1'h0;
    end else if (_T_3) begin
      if (io_en) begin
        if (startFlag) begin
          isDiv0 <= _T_4;
        end
      end
    end
    if (reset) begin
      lastDivident <= 32'h0;
    end else if (!(io_flush)) begin
      if (_T_3) begin
        if (io_en) begin
          if (startFlag) begin
            lastDivident <= io_divident;
          end
        end
      end
    end
    if (reset) begin
      lastDivisor <= 32'h0;
    end else if (!(io_flush)) begin
      if (_T_3) begin
        if (io_en) begin
          if (startFlag) begin
            lastDivisor <= io_divisor;
          end
        end
      end
    end
    if (reset) begin
      divisor <= 65'h0;
    end else if (!(io_flush)) begin
      if (_T_3) begin
        if (io_en) begin
          if (startFlag) begin
            if (!(_T_4)) begin
              divisor <= _T_8;
            end
          end
        end
      end
    end
  end
endmodule
module MDU(
  input         clock,
  input         reset,
  input         io_flush,
  input  [3:0]  io_op,
  output        io_valid,
  input  [31:0] io_opr1,
  input  [31:0] io_opr2,
  output [31:0] io_result
);
  wire  mul_clock; // @[MDU.scala 33:25]
  wire  mul_reset; // @[MDU.scala 33:25]
  wire  mul_io_en; // @[MDU.scala 33:25]
  wire  mul_io_flush; // @[MDU.scala 33:25]
  wire  mul_io_done; // @[MDU.scala 33:25]
  wire [31:0] mul_io_opr1; // @[MDU.scala 33:25]
  wire [31:0] mul_io_opr2; // @[MDU.scala 33:25]
  wire [63:0] mul_io_result; // @[MDU.scala 33:25]
  wire  div_clock; // @[MDU.scala 43:29]
  wire  div_reset; // @[MDU.scala 43:29]
  wire  div_io_en; // @[MDU.scala 43:29]
  wire  div_io_flush; // @[MDU.scala 43:29]
  wire  div_io_divZero; // @[MDU.scala 43:29]
  wire  div_io_done; // @[MDU.scala 43:29]
  wire [31:0] div_io_divident; // @[MDU.scala 43:29]
  wire [31:0] div_io_divisor; // @[MDU.scala 43:29]
  wire [31:0] div_io_quotient; // @[MDU.scala 43:29]
  wire [31:0] div_io_remainder; // @[MDU.scala 43:29]
  wire  _T_1 = 4'h1 == io_op; // @[Lookup.scala 31:38]
  wire  _T_3 = 4'h2 == io_op; // @[Lookup.scala 31:38]
  wire  _T_5 = 4'h3 == io_op; // @[Lookup.scala 31:38]
  wire  _T_7 = 4'h4 == io_op; // @[Lookup.scala 31:38]
  wire  _T_9 = 4'h5 == io_op; // @[Lookup.scala 31:38]
  wire  _T_11 = 4'h6 == io_op; // @[Lookup.scala 31:38]
  wire  _T_13 = 4'h7 == io_op; // @[Lookup.scala 31:38]
  wire  _T_15 = 4'h8 == io_op; // @[Lookup.scala 31:38]
  wire  _T_21 = _T_5 | _T_7; // @[Lookup.scala 33:37]
  wire  _T_22 = _T_3 | _T_21; // @[Lookup.scala 33:37]
  wire  mulEn = _T_1 | _T_22; // @[Lookup.scala 33:37]
  wire  _T_24 = _T_13 | _T_15; // @[Lookup.scala 33:37]
  wire  _T_25 = _T_11 | _T_24; // @[Lookup.scala 33:37]
  wire  _T_26 = _T_9 | _T_25; // @[Lookup.scala 33:37]
  wire  _T_27 = _T_7 ? 1'h0 : _T_26; // @[Lookup.scala 33:37]
  wire  _T_28 = _T_5 ? 1'h0 : _T_27; // @[Lookup.scala 33:37]
  wire  _T_29 = _T_3 ? 1'h0 : _T_28; // @[Lookup.scala 33:37]
  wire  divEn = _T_1 ? 1'h0 : _T_29; // @[Lookup.scala 33:37]
  wire  _T_32 = _T_11 ? 1'h0 : _T_24; // @[Lookup.scala 33:37]
  wire  _T_33 = _T_9 ? 1'h0 : _T_32; // @[Lookup.scala 33:37]
  wire  _T_34 = _T_7 | _T_33; // @[Lookup.scala 33:37]
  wire  _T_35 = _T_5 | _T_34; // @[Lookup.scala 33:37]
  wire  _T_36 = _T_3 | _T_35; // @[Lookup.scala 33:37]
  wire  hiRem = _T_1 ? 1'h0 : _T_36; // @[Lookup.scala 33:37]
  wire  _T_39 = _T_11 ? 1'h0 : _T_13; // @[Lookup.scala 33:37]
  wire  _T_40 = _T_9 | _T_39; // @[Lookup.scala 33:37]
  wire  _T_41 = _T_7 ? 1'h0 : _T_40; // @[Lookup.scala 33:37]
  wire  _T_42 = _T_5 | _T_41; // @[Lookup.scala 33:37]
  wire  _T_43 = _T_3 | _T_42; // @[Lookup.scala 33:37]
  wire  lhsSigned = _T_1 ? 1'h0 : _T_43; // @[Lookup.scala 33:37]
  wire  _T_49 = _T_5 ? 1'h0 : _T_41; // @[Lookup.scala 33:37]
  wire  _T_50 = _T_3 | _T_49; // @[Lookup.scala 33:37]
  wire  rhsSigned = _T_1 ? 1'h0 : _T_50; // @[Lookup.scala 33:37]
  wire  isOpr1Neg = lhsSigned & io_opr1[31]; // @[MDU.scala 26:29]
  wire  isOpr2Neg = rhsSigned & io_opr2[31]; // @[MDU.scala 27:29]
  wire  isAnsNeg = isOpr1Neg ^ isOpr2Neg; // @[MDU.scala 28:29]
  wire [31:0] _T_54 = 32'h0 - io_opr1; // @[MDU.scala 29:34]
  wire [31:0] opr1 = isOpr1Neg ? _T_54 : io_opr1; // @[MDU.scala 29:22]
  wire [31:0] _T_56 = 32'h0 - io_opr2; // @[MDU.scala 30:34]
  wire [31:0] opr2 = isOpr2Neg ? _T_56 : io_opr2; // @[MDU.scala 30:22]
  wire [63:0] _T_58 = 64'h0 - mul_io_result; // @[MDU.scala 34:33]
  wire [63:0] mulOut = isAnsNeg ? _T_58 : mul_io_result; // @[MDU.scala 34:22]
  wire [31:0] mulAns = hiRem ? mulOut[63:32] : mulOut[31:0]; // @[MDU.scala 35:22]
  wire  _T_61 = mulEn & mul_io_done; // @[MDU.scala 38:38]
  wire [32:0] _GEN_0 = {{1'd0}, opr1}; // @[MDU.scala 46:41]
  wire  _T_63 = _GEN_0 == 33'h100000000; // @[MDU.scala 46:41]
  wire  _T_64 = lhsSigned & _T_63; // @[MDU.scala 46:33]
  wire  _T_65 = opr2 == 32'hffffffff; // @[MDU.scala 46:60]
  wire  isDivOverflow = _T_64 & _T_65; // @[MDU.scala 46:52]
  wire  _T_68 = io_opr1[31] ^ div_io_remainder[31]; // @[MDU.scala 47:61]
  wire  isRemNeg = lhsSigned & _T_68; // @[MDU.scala 47:33]
  wire [31:0] _T_70 = 32'h0 - div_io_quotient; // @[MDU.scala 49:37]
  wire [31:0] divQuo = isAnsNeg ? _T_70 : div_io_quotient; // @[MDU.scala 49:26]
  wire [32:0] _T_71 = isDivOverflow ? 33'h100000000 : {{1'd0}, divQuo}; // @[MDU.scala 51:26]
  wire [32:0] divAnsQuo = div_io_divZero ? 33'hffffffff : _T_71; // @[MDU.scala 50:26]
  wire [31:0] _T_73 = 32'h0 - div_io_remainder; // @[MDU.scala 52:37]
  wire [31:0] divRem = isRemNeg ? _T_73 : div_io_remainder; // @[MDU.scala 52:26]
  wire [31:0] _T_74 = isDivOverflow ? 32'h0 : divRem; // @[MDU.scala 54:26]
  wire [31:0] divAnsRem = div_io_divZero ? io_opr1 : _T_74; // @[MDU.scala 53:26]
  wire [32:0] divAns = hiRem ? {{1'd0}, divAnsRem} : divAnsQuo; // @[MDU.scala 55:26]
  wire  _T_75 = divEn ? div_io_done : 1'h1; // @[MDU.scala 62:43]
  wire [32:0] _T_77 = divEn ? divAns : 33'h0; // @[MDU.scala 63:38]
  wire [32:0] _T_78 = mulEn ? {{1'd0}, mulAns} : _T_77; // @[MDU.scala 63:19]
  Multiplier mul ( // @[MDU.scala 33:25]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_en(mul_io_en),
    .io_flush(mul_io_flush),
    .io_done(mul_io_done),
    .io_opr1(mul_io_opr1),
    .io_opr2(mul_io_opr2),
    .io_result(mul_io_result)
  );
  Divider div ( // @[MDU.scala 43:29]
    .clock(div_clock),
    .reset(div_reset),
    .io_en(div_io_en),
    .io_flush(div_io_flush),
    .io_divZero(div_io_divZero),
    .io_done(div_io_done),
    .io_divident(div_io_divident),
    .io_divisor(div_io_divisor),
    .io_quotient(div_io_quotient),
    .io_remainder(div_io_remainder)
  );
  assign io_valid = mulEn ? mul_io_done : _T_75; // @[MDU.scala 62:13]
  assign io_result = _T_78[31:0]; // @[MDU.scala 63:13]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_en = _T_1 | _T_22; // @[MDU.scala 37:16]
  assign mul_io_flush = io_flush | _T_61; // @[MDU.scala 38:16]
  assign mul_io_opr1 = isOpr1Neg ? _T_54 : io_opr1; // @[MDU.scala 39:16]
  assign mul_io_opr2 = isOpr2Neg ? _T_56 : io_opr2; // @[MDU.scala 40:16]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_en = _T_1 ? 1'h0 : _T_29; // @[MDU.scala 56:20]
  assign div_io_flush = io_flush; // @[MDU.scala 57:20]
  assign div_io_divident = isOpr1Neg ? _T_54 : io_opr1; // @[MDU.scala 58:20]
  assign div_io_divisor = isOpr2Neg ? _T_56 : io_opr2; // @[MDU.scala 59:20]
endmodule
module ALU(
  input         clock,
  input         reset,
  input  [3:0]  io_decoder_aluOp,
  input  [31:0] io_decoder_opr1,
  input  [31:0] io_decoder_opr2,
  input  [3:0]  io_decoder_mduOp,
  input  [4:0]  io_decoder_lsuOp,
  input  [31:0] io_decoder_lsuData,
  input         io_decoder_regWen,
  input  [4:0]  io_decoder_regWaddr,
  input  [2:0]  io_decoder_csrOp,
  input  [11:0] io_decoder_csrAddr,
  input  [31:0] io_decoder_csrData,
  input  [3:0]  io_decoder_excType,
  input  [31:0] io_decoder_excValue,
  input         io_decoder_valid,
  input  [31:0] io_decoder_inst,
  input  [31:0] io_decoder_currentPc,
  input         io_flush,
  output        io_stallReq,
  output [2:0]  io_csrRead_op,
  input         io_csrRead_valid,
  output [11:0] io_csrRead_addr,
  input  [31:0] io_csrRead_data,
  output [4:0]  io_alu_lsuOp,
  output [31:0] io_alu_lsuData,
  output        io_alu_reg_en,
  output [4:0]  io_alu_reg_addr,
  output [31:0] io_alu_reg_data,
  output        io_alu_reg_load,
  output [2:0]  io_alu_csr_op,
  output [11:0] io_alu_csr_addr,
  output [31:0] io_alu_csr_data,
  output        io_alu_csr_retired,
  output [3:0]  io_alu_excType,
  output [31:0] io_alu_excValue,
  output        io_alu_valid,
  output [31:0] io_alu_inst,
  output [31:0] io_alu_currentPc
);
  wire  mdu_clock; // @[ALU.scala 48:25]
  wire  mdu_reset; // @[ALU.scala 48:25]
  wire  mdu_io_flush; // @[ALU.scala 48:25]
  wire [3:0] mdu_io_op; // @[ALU.scala 48:25]
  wire  mdu_io_valid; // @[ALU.scala 48:25]
  wire [31:0] mdu_io_opr1; // @[ALU.scala 48:25]
  wire [31:0] mdu_io_opr2; // @[ALU.scala 48:25]
  wire [31:0] mdu_io_result; // @[ALU.scala 48:25]
  wire [4:0] shamt = io_decoder_opr2[4:0]; // @[ALU.scala 31:19]
  wire [31:0] _T_1 = io_decoder_opr1 + io_decoder_opr2; // @[ALU.scala 35:24]
  wire [31:0] _T_3 = io_decoder_opr1 - io_decoder_opr2; // @[ALU.scala 36:24]
  wire [31:0] _T_4 = io_decoder_opr1 ^ io_decoder_opr2; // @[ALU.scala 37:24]
  wire [31:0] _T_5 = io_decoder_opr1 | io_decoder_opr2; // @[ALU.scala 38:24]
  wire [31:0] _T_6 = io_decoder_opr1 & io_decoder_opr2; // @[ALU.scala 39:24]
  wire  _T_9 = $signed(io_decoder_opr1) < $signed(io_decoder_opr2); // @[ALU.scala 40:31]
  wire  _T_10 = io_decoder_opr1 < io_decoder_opr2; // @[ALU.scala 41:24]
  wire [62:0] _GEN_0 = {{31'd0}, io_decoder_opr1}; // @[ALU.scala 42:24]
  wire [62:0] _T_11 = _GEN_0 << shamt; // @[ALU.scala 42:24]
  wire [31:0] _T_12 = io_decoder_opr1 >> shamt; // @[ALU.scala 43:24]
  wire [31:0] _T_15 = $signed(io_decoder_opr1) >>> shamt; // @[ALU.scala 44:41]
  wire  _T_16 = 4'h9 == io_decoder_aluOp; // @[Mux.scala 68:19]
  wire [31:0] _T_17 = _T_16 ? _T_15 : 32'h0; // @[Mux.scala 68:16]
  wire  _T_18 = 4'h8 == io_decoder_aluOp; // @[Mux.scala 68:19]
  wire [31:0] _T_19 = _T_18 ? _T_12 : _T_17; // @[Mux.scala 68:16]
  wire  _T_20 = 4'h7 == io_decoder_aluOp; // @[Mux.scala 68:19]
  wire [62:0] _T_21 = _T_20 ? _T_11 : {{31'd0}, _T_19}; // @[Mux.scala 68:16]
  wire  _T_22 = 4'h6 == io_decoder_aluOp; // @[Mux.scala 68:19]
  wire [62:0] _T_23 = _T_22 ? {{62'd0}, _T_10} : _T_21; // @[Mux.scala 68:16]
  wire  _T_24 = 4'h5 == io_decoder_aluOp; // @[Mux.scala 68:19]
  wire [62:0] _T_25 = _T_24 ? {{62'd0}, _T_9} : _T_23; // @[Mux.scala 68:16]
  wire  _T_26 = 4'h4 == io_decoder_aluOp; // @[Mux.scala 68:19]
  wire [62:0] _T_27 = _T_26 ? {{31'd0}, _T_6} : _T_25; // @[Mux.scala 68:16]
  wire  _T_28 = 4'h3 == io_decoder_aluOp; // @[Mux.scala 68:19]
  wire [62:0] _T_29 = _T_28 ? {{31'd0}, _T_5} : _T_27; // @[Mux.scala 68:16]
  wire  _T_30 = 4'h2 == io_decoder_aluOp; // @[Mux.scala 68:19]
  wire [62:0] _T_31 = _T_30 ? {{31'd0}, _T_4} : _T_29; // @[Mux.scala 68:16]
  wire  _T_32 = 4'h1 == io_decoder_aluOp; // @[Mux.scala 68:19]
  wire [62:0] _T_33 = _T_32 ? {{31'd0}, _T_3} : _T_31; // @[Mux.scala 68:16]
  wire  _T_34 = 4'h0 == io_decoder_aluOp; // @[Mux.scala 68:19]
  wire [62:0] aluResult = _T_34 ? {{31'd0}, _T_1} : _T_33; // @[Mux.scala 68:16]
  wire [31:0] mduResult = mdu_io_valid ? mdu_io_result : 32'h0; // @[ALU.scala 53:22]
  wire  csrEn = io_decoder_csrOp != 3'h0; // @[ALU.scala 56:34]
  wire  _T_35 = ~io_csrRead_valid; // @[ALU.scala 58:30]
  wire  _T_36 = csrEn & _T_35; // @[ALU.scala 58:27]
  wire  _T_37 = io_decoder_mduOp != 4'h0; // @[ALU.scala 63:38]
  wire [62:0] _T_38 = _T_37 ? {{31'd0}, mduResult} : aluResult; // @[ALU.scala 63:20]
  wire [62:0] result = csrEn ? {{31'd0}, io_csrRead_data} : _T_38; // @[ALU.scala 62:20]
  wire  _T_39 = io_decoder_lsuOp != 5'h0; // @[ALU.scala 64:34]
  MDU mdu ( // @[ALU.scala 48:25]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_flush(mdu_io_flush),
    .io_op(mdu_io_op),
    .io_valid(mdu_io_valid),
    .io_opr1(mdu_io_opr1),
    .io_opr2(mdu_io_opr2),
    .io_result(mdu_io_result)
  );
  assign io_stallReq = ~mdu_io_valid; // @[ALU.scala 67:15]
  assign io_csrRead_op = io_decoder_csrOp; // @[ALU.scala 70:19]
  assign io_csrRead_addr = io_decoder_csrAddr; // @[ALU.scala 71:19]
  assign io_alu_lsuOp = io_decoder_lsuOp; // @[ALU.scala 75:23]
  assign io_alu_lsuData = io_decoder_lsuData; // @[ALU.scala 76:23]
  assign io_alu_reg_en = io_decoder_regWen; // @[ALU.scala 78:23]
  assign io_alu_reg_addr = io_decoder_regWaddr; // @[ALU.scala 79:23]
  assign io_alu_reg_data = result[31:0]; // @[ALU.scala 80:23]
  assign io_alu_reg_load = _T_39 & io_decoder_regWen; // @[ALU.scala 81:23]
  assign io_alu_csr_op = io_decoder_csrOp; // @[ALU.scala 83:23]
  assign io_alu_csr_addr = io_decoder_csrAddr; // @[ALU.scala 84:23]
  assign io_alu_csr_data = io_decoder_csrData; // @[ALU.scala 85:23]
  assign io_alu_csr_retired = io_decoder_inst != 32'h13; // @[ALU.scala 86:23]
  assign io_alu_excType = _T_36 ? 4'h5 : io_decoder_excType; // @[ALU.scala 88:23]
  assign io_alu_excValue = io_decoder_excValue; // @[ALU.scala 89:23]
  assign io_alu_valid = io_decoder_valid; // @[ALU.scala 91:23]
  assign io_alu_inst = io_decoder_inst; // @[ALU.scala 92:23]
  assign io_alu_currentPc = io_decoder_currentPc; // @[ALU.scala 93:23]
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_flush = io_flush; // @[ALU.scala 49:17]
  assign mdu_io_op = io_decoder_mduOp; // @[ALU.scala 50:17]
  assign mdu_io_opr1 = io_decoder_opr1; // @[ALU.scala 51:17]
  assign mdu_io_opr2 = io_decoder_opr2; // @[ALU.scala 52:17]
endmodule
module MidStage_2(
  input         clock,
  input         reset,
  input         io_flush,
  input         io_stallPrev,
  input         io_stallNext,
  input  [4:0]  io_prev_lsuOp,
  input  [31:0] io_prev_lsuData,
  input         io_prev_reg_en,
  input  [4:0]  io_prev_reg_addr,
  input  [31:0] io_prev_reg_data,
  input  [2:0]  io_prev_csr_op,
  input  [11:0] io_prev_csr_addr,
  input  [31:0] io_prev_csr_data,
  input         io_prev_csr_retired,
  input  [3:0]  io_prev_excType,
  input  [31:0] io_prev_excValue,
  input         io_prev_valid,
  input  [31:0] io_prev_inst,
  input  [31:0] io_prev_currentPc,
  output [4:0]  io_next_lsuOp,
  output [31:0] io_next_lsuData,
  output        io_next_reg_en,
  output [4:0]  io_next_reg_addr,
  output [31:0] io_next_reg_data,
  output [2:0]  io_next_csr_op,
  output [11:0] io_next_csr_addr,
  output [31:0] io_next_csr_data,
  output        io_next_csr_retired,
  output [3:0]  io_next_excType,
  output [31:0] io_next_excValue,
  output        io_next_valid,
  output [31:0] io_next_inst,
  output [31:0] io_next_currentPc
);
  reg [4:0] ff_lsuOp; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_0;
  reg [31:0] ff_lsuData; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_1;
  reg  ff_reg_en; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_2;
  reg [4:0] ff_reg_addr; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_3;
  reg [31:0] ff_reg_data; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_4;
  reg [2:0] ff_csr_op; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_5;
  reg [11:0] ff_csr_addr; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_6;
  reg [31:0] ff_csr_data; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_7;
  reg  ff_csr_retired; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_8;
  reg [3:0] ff_excType; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_9;
  reg [31:0] ff_excValue; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_10;
  reg  ff_valid; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_11;
  reg [31:0] ff_inst; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_12;
  reg [31:0] ff_currentPc; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_13;
  wire  _T_1 = ~io_stallNext; // @[MidStage.scala 21:38]
  wire  _T_2 = io_stallPrev & _T_1; // @[MidStage.scala 21:35]
  wire  _T_3 = io_flush | _T_2; // @[MidStage.scala 21:18]
  wire  _T_5 = ~io_stallPrev; // @[MidStage.scala 23:15]
  assign io_next_lsuOp = ff_lsuOp; // @[MidStage.scala 27:11]
  assign io_next_lsuData = ff_lsuData; // @[MidStage.scala 27:11]
  assign io_next_reg_en = ff_reg_en; // @[MidStage.scala 27:11]
  assign io_next_reg_addr = ff_reg_addr; // @[MidStage.scala 27:11]
  assign io_next_reg_data = ff_reg_data; // @[MidStage.scala 27:11]
  assign io_next_csr_op = ff_csr_op; // @[MidStage.scala 27:11]
  assign io_next_csr_addr = ff_csr_addr; // @[MidStage.scala 27:11]
  assign io_next_csr_data = ff_csr_data; // @[MidStage.scala 27:11]
  assign io_next_csr_retired = ff_csr_retired; // @[MidStage.scala 27:11]
  assign io_next_excType = ff_excType; // @[MidStage.scala 27:11]
  assign io_next_excValue = ff_excValue; // @[MidStage.scala 27:11]
  assign io_next_valid = ff_valid; // @[MidStage.scala 27:11]
  assign io_next_inst = ff_inst; // @[MidStage.scala 27:11]
  assign io_next_currentPc = ff_currentPc; // @[MidStage.scala 27:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff_lsuOp = _RAND_0[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ff_lsuData = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ff_reg_en = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ff_reg_addr = _RAND_3[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ff_reg_data = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ff_csr_op = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ff_csr_addr = _RAND_6[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ff_csr_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ff_csr_retired = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  ff_excType = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  ff_excValue = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  ff_valid = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  ff_inst = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  ff_currentPc = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ff_lsuOp <= 5'h0;
    end else if (_T_3) begin
      ff_lsuOp <= 5'h0;
    end else if (_T_5) begin
      ff_lsuOp <= io_prev_lsuOp;
    end
    if (reset) begin
      ff_lsuData <= 32'h0;
    end else if (_T_3) begin
      ff_lsuData <= 32'h0;
    end else if (_T_5) begin
      ff_lsuData <= io_prev_lsuData;
    end
    if (reset) begin
      ff_reg_en <= 1'h0;
    end else if (_T_3) begin
      ff_reg_en <= 1'h0;
    end else if (_T_5) begin
      ff_reg_en <= io_prev_reg_en;
    end
    if (reset) begin
      ff_reg_addr <= 5'h0;
    end else if (_T_3) begin
      ff_reg_addr <= 5'h0;
    end else if (_T_5) begin
      ff_reg_addr <= io_prev_reg_addr;
    end
    if (reset) begin
      ff_reg_data <= 32'h0;
    end else if (_T_3) begin
      ff_reg_data <= 32'h0;
    end else if (_T_5) begin
      ff_reg_data <= io_prev_reg_data;
    end
    if (reset) begin
      ff_csr_op <= 3'h0;
    end else if (_T_3) begin
      ff_csr_op <= 3'h0;
    end else if (_T_5) begin
      ff_csr_op <= io_prev_csr_op;
    end
    if (reset) begin
      ff_csr_addr <= 12'h0;
    end else if (_T_3) begin
      ff_csr_addr <= 12'h0;
    end else if (_T_5) begin
      ff_csr_addr <= io_prev_csr_addr;
    end
    if (reset) begin
      ff_csr_data <= 32'h0;
    end else if (_T_3) begin
      ff_csr_data <= 32'h0;
    end else if (_T_5) begin
      ff_csr_data <= io_prev_csr_data;
    end
    if (reset) begin
      ff_csr_retired <= 1'h0;
    end else if (_T_3) begin
      ff_csr_retired <= 1'h0;
    end else if (_T_5) begin
      ff_csr_retired <= io_prev_csr_retired;
    end
    if (reset) begin
      ff_excType <= 4'h0;
    end else if (_T_3) begin
      ff_excType <= 4'h0;
    end else if (_T_5) begin
      ff_excType <= io_prev_excType;
    end
    if (reset) begin
      ff_excValue <= 32'h0;
    end else if (_T_3) begin
      ff_excValue <= 32'h0;
    end else if (_T_5) begin
      ff_excValue <= io_prev_excValue;
    end
    if (reset) begin
      ff_valid <= 1'h0;
    end else if (_T_3) begin
      ff_valid <= 1'h0;
    end else if (_T_5) begin
      ff_valid <= io_prev_valid;
    end
    if (reset) begin
      ff_inst <= 32'h0;
    end else if (_T_3) begin
      ff_inst <= 32'h0;
    end else if (_T_5) begin
      ff_inst <= io_prev_inst;
    end
    if (reset) begin
      ff_currentPc <= 32'h0;
    end else if (_T_3) begin
      ff_currentPc <= 32'h0;
    end else if (_T_5) begin
      ff_currentPc <= io_prev_currentPc;
    end
  end
endmodule
module AmoExecute(
  input         clock,
  input         reset,
  input  [3:0]  io_op,
  input         io_flush,
  output        io_ready,
  input  [31:0] io_regOpr,
  output [31:0] io_regWdata,
  input         io_ramValid,
  output        io_ramWen,
  input  [31:0] io_ramRdata,
  output [31:0] io_ramWdata
);
  reg [1:0] state; // @[AmoExecute.scala 28:22]
  reg [31:0] _RAND_0;
  wire [31:0] _T_1 = io_ramRdata + io_regOpr; // @[AmoExecute.scala 37:26]
  wire [31:0] _T_2 = io_ramRdata ^ io_regOpr; // @[AmoExecute.scala 38:26]
  wire [31:0] _T_3 = io_ramRdata & io_regOpr; // @[AmoExecute.scala 39:26]
  wire [31:0] _T_4 = io_ramRdata | io_regOpr; // @[AmoExecute.scala 40:26]
  wire  _T_7 = $signed(io_ramRdata) < $signed(io_regOpr); // @[AmoExecute.scala 41:36]
  wire [31:0] _T_8 = _T_7 ? io_ramRdata : io_regOpr; // @[AmoExecute.scala 41:23]
  wire  _T_11 = $signed(io_ramRdata) > $signed(io_regOpr); // @[AmoExecute.scala 42:36]
  wire [31:0] _T_12 = _T_11 ? io_ramRdata : io_regOpr; // @[AmoExecute.scala 42:23]
  wire  _T_13 = io_ramRdata < io_regOpr; // @[AmoExecute.scala 43:29]
  wire [31:0] _T_14 = _T_13 ? io_ramRdata : io_regOpr; // @[AmoExecute.scala 43:23]
  wire  _T_15 = io_ramRdata > io_regOpr; // @[AmoExecute.scala 44:29]
  wire [31:0] _T_16 = _T_15 ? io_ramRdata : io_regOpr; // @[AmoExecute.scala 44:23]
  wire  _T_17 = 4'h9 == io_op; // @[Mux.scala 68:19]
  wire [31:0] _T_18 = _T_17 ? _T_16 : 32'h0; // @[Mux.scala 68:16]
  wire  _T_19 = 4'h8 == io_op; // @[Mux.scala 68:19]
  wire [31:0] _T_20 = _T_19 ? _T_14 : _T_18; // @[Mux.scala 68:16]
  wire  _T_21 = 4'h7 == io_op; // @[Mux.scala 68:19]
  wire [31:0] _T_22 = _T_21 ? _T_12 : _T_20; // @[Mux.scala 68:16]
  wire  _T_23 = 4'h6 == io_op; // @[Mux.scala 68:19]
  wire [31:0] _T_24 = _T_23 ? _T_8 : _T_22; // @[Mux.scala 68:16]
  wire  _T_25 = 4'h5 == io_op; // @[Mux.scala 68:19]
  wire [31:0] _T_26 = _T_25 ? _T_4 : _T_24; // @[Mux.scala 68:16]
  wire  _T_27 = 4'h4 == io_op; // @[Mux.scala 68:19]
  wire [31:0] _T_28 = _T_27 ? _T_3 : _T_26; // @[Mux.scala 68:16]
  wire  _T_29 = 4'h3 == io_op; // @[Mux.scala 68:19]
  wire [31:0] _T_30 = _T_29 ? _T_2 : _T_28; // @[Mux.scala 68:16]
  wire  _T_31 = 4'h2 == io_op; // @[Mux.scala 68:19]
  wire [31:0] _T_32 = _T_31 ? _T_1 : _T_30; // @[Mux.scala 68:16]
  wire  _T_33 = 4'h1 == io_op; // @[Mux.scala 68:19]
  wire  _T_34 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_35 = io_op == 4'h0; // @[AmoExecute.scala 56:21]
  wire  _T_36 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_37 = 2'h2 == state; // @[Conditional.scala 37:30]
  assign io_ready = state == 2'h2; // @[AmoExecute.scala 75:15]
  assign io_regWdata = io_ramRdata; // @[AmoExecute.scala 76:15]
  assign io_ramWen = state == 2'h1; // @[AmoExecute.scala 77:15]
  assign io_ramWdata = _T_33 ? io_regOpr : _T_32; // @[AmoExecute.scala 78:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (io_flush) begin
      state <= 2'h0;
    end else if (io_ramValid) begin
      if (_T_34) begin
        if (_T_35) begin
          state <= 2'h0;
        end else begin
          state <= 2'h1;
        end
      end else if (_T_36) begin
        state <= 2'h2;
      end else if (_T_37) begin
        state <= 2'h0;
      end
    end
  end
endmodule
module Mem(
  input         clock,
  input         reset,
  input  [4:0]  io_alu_lsuOp,
  input  [31:0] io_alu_lsuData,
  input         io_alu_reg_en,
  input  [4:0]  io_alu_reg_addr,
  input  [31:0] io_alu_reg_data,
  input  [2:0]  io_alu_csr_op,
  input  [11:0] io_alu_csr_addr,
  input  [31:0] io_alu_csr_data,
  input         io_alu_csr_retired,
  input  [3:0]  io_alu_excType,
  input  [31:0] io_alu_excValue,
  input         io_alu_valid,
  input  [31:0] io_alu_inst,
  input  [31:0] io_alu_currentPc,
  input         io_flush,
  output        io_stallReq,
  output        io_flushReq,
  output [31:0] io_flushPc,
  output        io_ram_en,
  input         io_ram_valid,
  input         io_ram_fault,
  output [3:0]  io_ram_wen,
  output [31:0] io_ram_addr,
  input  [31:0] io_ram_rdata,
  output [31:0] io_ram_wdata,
  output        io_flushIc,
  output        io_flushDc,
  output        io_flushIt,
  output        io_flushDt,
  input         io_csrHasInt,
  input         io_csrBusy,
  input  [1:0]  io_csrMode,
  output [31:0] io_excMon_addr,
  input         io_excMon_valid,
  output        io_except_hasTrap,
  output        io_except_isSret,
  output        io_except_isMret,
  output [30:0] io_except_excCause,
  output [31:0] io_except_excPc,
  output [31:0] io_except_excValue,
  output        io_mem_reg_en,
  output [4:0]  io_mem_reg_addr,
  output [31:0] io_mem_reg_data,
  output        io_mem_reg_load,
  output        io_mem_memSigned,
  output [1:0]  io_mem_memSel,
  output [1:0]  io_mem_memWidth,
  output [2:0]  io_mem_csr_op,
  output [11:0] io_mem_csr_addr,
  output [31:0] io_mem_csr_data,
  output        io_mem_csr_retired,
  output [31:0] io_mem_excMon_addr,
  output        io_mem_excMon_set,
  output        io_mem_excMon_clear,
  output [31:0] io_mem_currentPc
);
  wire  amo_clock; // @[Mem.scala 55:19]
  wire  amo_reset; // @[Mem.scala 55:19]
  wire [3:0] amo_io_op; // @[Mem.scala 55:19]
  wire  amo_io_flush; // @[Mem.scala 55:19]
  wire  amo_io_ready; // @[Mem.scala 55:19]
  wire [31:0] amo_io_regOpr; // @[Mem.scala 55:19]
  wire [31:0] amo_io_regWdata; // @[Mem.scala 55:19]
  wire  amo_io_ramValid; // @[Mem.scala 55:19]
  wire  amo_io_ramWen; // @[Mem.scala 55:19]
  wire [31:0] amo_io_ramRdata; // @[Mem.scala 55:19]
  wire [31:0] amo_io_ramWdata; // @[Mem.scala 55:19]
  wire  _T_1 = 5'h1 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_3 = 5'h2 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_5 = 5'h3 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_7 = 5'h4 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_9 = 5'h5 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_11 = 5'h6 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_13 = 5'h7 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_15 = 5'h8 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_17 = 5'h9 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_19 = 5'ha == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_21 = 5'hb == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_23 = 5'hc == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_25 = 5'hd == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_27 = 5'he == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_29 = 5'hf == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_31 = 5'h10 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_33 = 5'h11 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_35 = 5'h12 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_37 = 5'h13 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_39 = 5'h14 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_41 = 5'h15 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_43 = 5'h16 == io_alu_lsuOp; // @[Lookup.scala 31:38]
  wire  _T_48 = _T_35 | _T_37; // @[Lookup.scala 33:37]
  wire  _T_49 = _T_33 | _T_48; // @[Lookup.scala 33:37]
  wire  _T_50 = _T_31 | _T_49; // @[Lookup.scala 33:37]
  wire  _T_51 = _T_29 | _T_50; // @[Lookup.scala 33:37]
  wire  _T_52 = _T_27 | _T_51; // @[Lookup.scala 33:37]
  wire  _T_53 = _T_25 | _T_52; // @[Lookup.scala 33:37]
  wire  _T_54 = _T_23 | _T_53; // @[Lookup.scala 33:37]
  wire  _T_55 = _T_21 | _T_54; // @[Lookup.scala 33:37]
  wire  _T_56 = _T_19 | _T_55; // @[Lookup.scala 33:37]
  wire  _T_57 = _T_17 | _T_56; // @[Lookup.scala 33:37]
  wire  _T_58 = _T_15 | _T_57; // @[Lookup.scala 33:37]
  wire  _T_59 = _T_13 | _T_58; // @[Lookup.scala 33:37]
  wire  _T_60 = _T_11 | _T_59; // @[Lookup.scala 33:37]
  wire  _T_61 = _T_9 | _T_60; // @[Lookup.scala 33:37]
  wire  _T_62 = _T_7 | _T_61; // @[Lookup.scala 33:37]
  wire  _T_63 = _T_5 | _T_62; // @[Lookup.scala 33:37]
  wire  _T_64 = _T_3 | _T_63; // @[Lookup.scala 33:37]
  wire  en = _T_1 | _T_64; // @[Lookup.scala 33:37]
  wire  _T_80 = _T_13 | _T_15; // @[Lookup.scala 33:37]
  wire  _T_81 = _T_11 | _T_80; // @[Lookup.scala 33:37]
  wire  _T_82 = _T_9 ? 1'h0 : _T_81; // @[Lookup.scala 33:37]
  wire  _T_83 = _T_7 ? 1'h0 : _T_82; // @[Lookup.scala 33:37]
  wire  _T_84 = _T_5 ? 1'h0 : _T_83; // @[Lookup.scala 33:37]
  wire  _T_85 = _T_3 ? 1'h0 : _T_84; // @[Lookup.scala 33:37]
  wire  wen = _T_1 ? 1'h0 : _T_85; // @[Lookup.scala 33:37]
  wire  _T_100 = _T_15 ? 1'h0 : _T_17; // @[Lookup.scala 33:37]
  wire  _T_101 = _T_13 ? 1'h0 : _T_100; // @[Lookup.scala 33:37]
  wire  _T_102 = _T_11 ? 1'h0 : _T_101; // @[Lookup.scala 33:37]
  wire  _T_103 = _T_9 | _T_102; // @[Lookup.scala 33:37]
  wire  _T_104 = _T_7 | _T_103; // @[Lookup.scala 33:37]
  wire  _T_105 = _T_5 | _T_104; // @[Lookup.scala 33:37]
  wire  _T_106 = _T_3 | _T_105; // @[Lookup.scala 33:37]
  wire [1:0] _T_110 = _T_37 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _T_111 = _T_35 ? 2'h2 : _T_110; // @[Lookup.scala 33:37]
  wire [1:0] _T_112 = _T_33 ? 2'h2 : _T_111; // @[Lookup.scala 33:37]
  wire [1:0] _T_113 = _T_31 ? 2'h2 : _T_112; // @[Lookup.scala 33:37]
  wire [1:0] _T_114 = _T_29 ? 2'h2 : _T_113; // @[Lookup.scala 33:37]
  wire [1:0] _T_115 = _T_27 ? 2'h2 : _T_114; // @[Lookup.scala 33:37]
  wire [1:0] _T_116 = _T_25 ? 2'h2 : _T_115; // @[Lookup.scala 33:37]
  wire [1:0] _T_117 = _T_23 ? 2'h2 : _T_116; // @[Lookup.scala 33:37]
  wire [1:0] _T_118 = _T_21 ? 2'h2 : _T_117; // @[Lookup.scala 33:37]
  wire [1:0] _T_119 = _T_19 ? 2'h2 : _T_118; // @[Lookup.scala 33:37]
  wire [1:0] _T_120 = _T_17 ? 2'h2 : _T_119; // @[Lookup.scala 33:37]
  wire [1:0] _T_121 = _T_15 ? 2'h2 : _T_120; // @[Lookup.scala 33:37]
  wire [1:0] _T_122 = _T_13 ? 2'h1 : _T_121; // @[Lookup.scala 33:37]
  wire [1:0] _T_123 = _T_11 ? 2'h0 : _T_122; // @[Lookup.scala 33:37]
  wire [1:0] _T_124 = _T_9 ? 2'h1 : _T_123; // @[Lookup.scala 33:37]
  wire [1:0] _T_125 = _T_7 ? 2'h0 : _T_124; // @[Lookup.scala 33:37]
  wire [1:0] _T_126 = _T_5 ? 2'h2 : _T_125; // @[Lookup.scala 33:37]
  wire [1:0] _T_127 = _T_3 ? 2'h1 : _T_126; // @[Lookup.scala 33:37]
  wire [1:0] width = _T_1 ? 2'h0 : _T_127; // @[Lookup.scala 33:37]
  wire  _T_166 = _T_9 ? 1'h0 : _T_102; // @[Lookup.scala 33:37]
  wire  _T_167 = _T_7 ? 1'h0 : _T_166; // @[Lookup.scala 33:37]
  wire  _T_168 = _T_5 ? 1'h0 : _T_167; // @[Lookup.scala 33:37]
  wire  _T_169 = _T_3 ? 1'h0 : _T_168; // @[Lookup.scala 33:37]
  wire  _T_183 = _T_17 ? 1'h0 : _T_19; // @[Lookup.scala 33:37]
  wire  _T_184 = _T_15 ? 1'h0 : _T_183; // @[Lookup.scala 33:37]
  wire  _T_185 = _T_13 ? 1'h0 : _T_184; // @[Lookup.scala 33:37]
  wire  _T_186 = _T_11 ? 1'h0 : _T_185; // @[Lookup.scala 33:37]
  wire  _T_187 = _T_9 ? 1'h0 : _T_186; // @[Lookup.scala 33:37]
  wire  _T_188 = _T_7 ? 1'h0 : _T_187; // @[Lookup.scala 33:37]
  wire  _T_189 = _T_5 ? 1'h0 : _T_188; // @[Lookup.scala 33:37]
  wire  _T_190 = _T_3 ? 1'h0 : _T_189; // @[Lookup.scala 33:37]
  wire  checkExcMon = _T_1 ? 1'h0 : _T_190; // @[Lookup.scala 33:37]
  wire [3:0] _T_194 = _T_37 ? 4'h9 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_195 = _T_35 ? 4'h8 : _T_194; // @[Lookup.scala 33:37]
  wire [3:0] _T_196 = _T_33 ? 4'h7 : _T_195; // @[Lookup.scala 33:37]
  wire [3:0] _T_197 = _T_31 ? 4'h6 : _T_196; // @[Lookup.scala 33:37]
  wire [3:0] _T_198 = _T_29 ? 4'h5 : _T_197; // @[Lookup.scala 33:37]
  wire [3:0] _T_199 = _T_27 ? 4'h4 : _T_198; // @[Lookup.scala 33:37]
  wire [3:0] _T_200 = _T_25 ? 4'h3 : _T_199; // @[Lookup.scala 33:37]
  wire [3:0] _T_201 = _T_23 ? 4'h2 : _T_200; // @[Lookup.scala 33:37]
  wire [3:0] _T_202 = _T_21 ? 4'h1 : _T_201; // @[Lookup.scala 33:37]
  wire [3:0] _T_203 = _T_19 ? 4'h0 : _T_202; // @[Lookup.scala 33:37]
  wire [3:0] _T_204 = _T_17 ? 4'h0 : _T_203; // @[Lookup.scala 33:37]
  wire [3:0] _T_205 = _T_15 ? 4'h0 : _T_204; // @[Lookup.scala 33:37]
  wire [3:0] _T_206 = _T_13 ? 4'h0 : _T_205; // @[Lookup.scala 33:37]
  wire [3:0] _T_207 = _T_11 ? 4'h0 : _T_206; // @[Lookup.scala 33:37]
  wire [3:0] _T_208 = _T_9 ? 4'h0 : _T_207; // @[Lookup.scala 33:37]
  wire [3:0] _T_209 = _T_7 ? 4'h0 : _T_208; // @[Lookup.scala 33:37]
  wire [3:0] _T_210 = _T_5 ? 4'h0 : _T_209; // @[Lookup.scala 33:37]
  wire [3:0] _T_211 = _T_3 ? 4'h0 : _T_210; // @[Lookup.scala 33:37]
  wire [3:0] amoOp = _T_1 ? 4'h0 : _T_211; // @[Lookup.scala 33:37]
  wire  _T_213 = _T_41 | _T_43; // @[Lookup.scala 33:37]
  wire  _T_214 = _T_39 ? 1'h0 : _T_213; // @[Lookup.scala 33:37]
  wire  _T_215 = _T_37 ? 1'h0 : _T_214; // @[Lookup.scala 33:37]
  wire  _T_216 = _T_35 ? 1'h0 : _T_215; // @[Lookup.scala 33:37]
  wire  _T_217 = _T_33 ? 1'h0 : _T_216; // @[Lookup.scala 33:37]
  wire  _T_218 = _T_31 ? 1'h0 : _T_217; // @[Lookup.scala 33:37]
  wire  _T_219 = _T_29 ? 1'h0 : _T_218; // @[Lookup.scala 33:37]
  wire  _T_220 = _T_27 ? 1'h0 : _T_219; // @[Lookup.scala 33:37]
  wire  _T_221 = _T_25 ? 1'h0 : _T_220; // @[Lookup.scala 33:37]
  wire  _T_222 = _T_23 ? 1'h0 : _T_221; // @[Lookup.scala 33:37]
  wire  _T_223 = _T_21 ? 1'h0 : _T_222; // @[Lookup.scala 33:37]
  wire  _T_224 = _T_19 ? 1'h0 : _T_223; // @[Lookup.scala 33:37]
  wire  _T_225 = _T_17 ? 1'h0 : _T_224; // @[Lookup.scala 33:37]
  wire  _T_226 = _T_15 ? 1'h0 : _T_225; // @[Lookup.scala 33:37]
  wire  _T_227 = _T_13 ? 1'h0 : _T_226; // @[Lookup.scala 33:37]
  wire  _T_228 = _T_11 ? 1'h0 : _T_227; // @[Lookup.scala 33:37]
  wire  _T_229 = _T_9 ? 1'h0 : _T_228; // @[Lookup.scala 33:37]
  wire  _T_230 = _T_7 ? 1'h0 : _T_229; // @[Lookup.scala 33:37]
  wire  _T_231 = _T_5 ? 1'h0 : _T_230; // @[Lookup.scala 33:37]
  wire  _T_232 = _T_3 ? 1'h0 : _T_231; // @[Lookup.scala 33:37]
  wire  flushIc = _T_1 ? 1'h0 : _T_232; // @[Lookup.scala 33:37]
  wire  _T_255 = _T_41 ? 1'h0 : _T_43; // @[Lookup.scala 33:37]
  wire  _T_256 = _T_39 ? 1'h0 : _T_255; // @[Lookup.scala 33:37]
  wire  _T_257 = _T_37 ? 1'h0 : _T_256; // @[Lookup.scala 33:37]
  wire  _T_258 = _T_35 ? 1'h0 : _T_257; // @[Lookup.scala 33:37]
  wire  _T_259 = _T_33 ? 1'h0 : _T_258; // @[Lookup.scala 33:37]
  wire  _T_260 = _T_31 ? 1'h0 : _T_259; // @[Lookup.scala 33:37]
  wire  _T_261 = _T_29 ? 1'h0 : _T_260; // @[Lookup.scala 33:37]
  wire  _T_262 = _T_27 ? 1'h0 : _T_261; // @[Lookup.scala 33:37]
  wire  _T_263 = _T_25 ? 1'h0 : _T_262; // @[Lookup.scala 33:37]
  wire  _T_264 = _T_23 ? 1'h0 : _T_263; // @[Lookup.scala 33:37]
  wire  _T_265 = _T_21 ? 1'h0 : _T_264; // @[Lookup.scala 33:37]
  wire  _T_266 = _T_19 ? 1'h0 : _T_265; // @[Lookup.scala 33:37]
  wire  _T_267 = _T_17 ? 1'h0 : _T_266; // @[Lookup.scala 33:37]
  wire  _T_268 = _T_15 ? 1'h0 : _T_267; // @[Lookup.scala 33:37]
  wire  _T_269 = _T_13 ? 1'h0 : _T_268; // @[Lookup.scala 33:37]
  wire  _T_270 = _T_11 ? 1'h0 : _T_269; // @[Lookup.scala 33:37]
  wire  _T_271 = _T_9 ? 1'h0 : _T_270; // @[Lookup.scala 33:37]
  wire  _T_272 = _T_7 ? 1'h0 : _T_271; // @[Lookup.scala 33:37]
  wire  _T_273 = _T_5 ? 1'h0 : _T_272; // @[Lookup.scala 33:37]
  wire  _T_274 = _T_3 ? 1'h0 : _T_273; // @[Lookup.scala 33:37]
  wire  flushIt = _T_1 ? 1'h0 : _T_274; // @[Lookup.scala 33:37]
  wire [1:0] sel = io_alu_reg_data[1:0]; // @[Mem.scala 52:30]
  wire [6:0] _T_297 = 7'h1 << sel; // @[Mem.scala 65:49]
  wire [6:0] _T_298 = 7'h3 << sel; // @[Mem.scala 66:50]
  wire  _T_299 = 2'h2 == width; // @[Mux.scala 68:19]
  wire [3:0] _T_300 = _T_299 ? 4'hf : 4'h0; // @[Mux.scala 68:16]
  wire  _T_301 = 2'h1 == width; // @[Mux.scala 68:19]
  wire [6:0] _T_302 = _T_301 ? _T_298 : {{3'd0}, _T_300}; // @[Mux.scala 68:16]
  wire  _T_303 = 2'h0 == width; // @[Mux.scala 68:19]
  wire [6:0] writeEn = _T_303 ? _T_297 : _T_302; // @[Mux.scala 68:16]
  wire [3:0] scWen = io_excMon_valid ? 4'hf : 4'h0; // @[Mem.scala 69:20]
  wire [3:0] amoWen = amo_io_ramWen ? 4'hf : 4'h0; // @[Mem.scala 70:20]
  wire [3:0] _T_304 = checkExcMon ? scWen : amoWen; // @[Mem.scala 71:38]
  wire [6:0] ramWen = wen ? writeEn : {{3'd0}, _T_304}; // @[Mem.scala 71:20]
  wire [39:0] _T_306 = {io_alu_lsuData, 8'h0}; // @[Mem.scala 75:40]
  wire [47:0] _T_307 = {io_alu_lsuData, 16'h0}; // @[Mem.scala 75:40]
  wire [55:0] _T_308 = {io_alu_lsuData, 24'h0}; // @[Mem.scala 75:40]
  wire  _T_312 = 2'h3 == sel; // @[Mux.scala 68:19]
  wire [55:0] _T_313 = _T_312 ? _T_308 : 56'h0; // @[Mux.scala 68:16]
  wire  _T_314 = 2'h2 == sel; // @[Mux.scala 68:19]
  wire [55:0] _T_315 = _T_314 ? {{8'd0}, _T_307} : _T_313; // @[Mux.scala 68:16]
  wire  _T_316 = 2'h1 == sel; // @[Mux.scala 68:19]
  wire [55:0] _T_317 = _T_316 ? {{16'd0}, _T_306} : _T_315; // @[Mux.scala 68:16]
  wire  _T_318 = 2'h0 == sel; // @[Mux.scala 68:19]
  wire [55:0] _T_319 = _T_318 ? {{24'd0}, io_alu_lsuData} : _T_317; // @[Mux.scala 68:16]
  wire [47:0] _T_321 = _T_314 ? _T_307 : 48'h0; // @[Mux.scala 68:16]
  wire [47:0] _T_323 = _T_318 ? {{16'd0}, io_alu_lsuData} : _T_321; // @[Mux.scala 68:16]
  wire [31:0] _T_325 = _T_318 ? io_alu_lsuData : 32'h0; // @[Mux.scala 68:16]
  wire [31:0] _T_327 = _T_299 ? _T_325 : 32'h0; // @[Mux.scala 68:16]
  wire [47:0] _T_329 = _T_301 ? _T_323 : {{16'd0}, _T_327}; // @[Mux.scala 68:16]
  wire [55:0] lsuData = _T_303 ? _T_319 : {{8'd0}, _T_329}; // @[Mux.scala 68:16]
  wire  _T_331 = wen | checkExcMon; // @[Mem.scala 84:25]
  wire [55:0] wdata = _T_331 ? lsuData : {{24'd0}, amo_io_ramWdata}; // @[Mem.scala 84:20]
  wire  _T_332 = amoOp != 4'h0; // @[Mem.scala 87:29]
  wire  _T_333 = ~amo_io_ready; // @[Mem.scala 87:45]
  wire  _T_334 = ~io_ram_valid; // @[Mem.scala 88:29]
  wire  _T_335 = en & _T_334; // @[Mem.scala 88:26]
  wire  memStall = _T_332 ? _T_333 : _T_335; // @[Mem.scala 87:22]
  wire  fencStall = flushIc & _T_334; // @[Mem.scala 89:27]
  wire  _T_337 = memStall | fencStall; // @[Mem.scala 90:28]
  wire  stallReq = _T_337 | io_csrBusy; // @[Mem.scala 90:41]
  wire  _T_338 = io_excMon_valid ? 1'h0 : 1'h1; // @[Mem.scala 93:34]
  wire [31:0] _T_340 = _T_332 ? amo_io_regWdata : io_alu_reg_data; // @[Mem.scala 94:17]
  wire  _T_346 = sel != 2'h0; // @[Mem.scala 104:33]
  wire  _T_348 = _T_299 & _T_346; // @[Mux.scala 68:16]
  wire  _T_350 = _T_301 ? sel[0] : _T_348; // @[Mux.scala 68:16]
  wire  memAddr = _T_303 ? 1'h0 : _T_350; // @[Mux.scala 68:16]
  wire  memExcept = memAddr | io_ram_fault; // @[Mem.scala 106:27]
  wire  _T_352 = io_alu_excType == 4'h3; // @[Mem.scala 108:34]
  wire  _T_353 = io_csrMode == 2'h0; // @[Mem.scala 108:61]
  wire  illgSret = _T_352 & _T_353; // @[Mem.scala 108:47]
  wire  _T_354 = io_alu_excType == 4'h4; // @[Mem.scala 109:34]
  wire  _T_355 = io_csrMode != 2'h3; // @[Mem.scala 109:61]
  wire  illgMret = _T_354 & _T_355; // @[Mem.scala 109:47]
  wire  _T_356 = io_alu_excType == 4'ha; // @[Mem.scala 110:34]
  wire  illgSpriv = _T_356 & _T_353; // @[Mem.scala 110:48]
  wire  instAddr = io_alu_excType == 4'h7; // @[Mem.scala 111:34]
  wire  instPage = io_alu_excType == 4'h6; // @[Mem.scala 112:34]
  wire  _T_358 = io_alu_excType == 4'h5; // @[Mem.scala 113:34]
  wire  _T_359 = _T_358 | illgSret; // @[Mem.scala 113:48]
  wire  _T_360 = _T_359 | illgMret; // @[Mem.scala 114:28]
  wire  instIllg = _T_360 | illgSpriv; // @[Mem.scala 114:40]
  wire  _T_361 = io_alu_excType == 4'h8; // @[Mem.scala 116:34]
  wire  _T_362 = io_alu_excType == 4'h9; // @[Mem.scala 117:34]
  wire  excMem = _T_361 | _T_362; // @[Mem.scala 116:47]
  wire  _T_363 = io_alu_excType == 4'h1; // @[Mem.scala 118:34]
  wire  _T_364 = io_alu_excType == 4'h2; // @[Mem.scala 119:34]
  wire  _T_365 = _T_363 | _T_364; // @[Mem.scala 118:48]
  wire  _T_367 = _T_365 | _T_352; // @[Mem.scala 119:47]
  wire  excOther = _T_367 | _T_354; // @[Mem.scala 120:47]
  wire  _T_369 = instAddr | instIllg; // @[Mem.scala 122:28]
  wire  _T_370 = _T_369 | instPage; // @[Mem.scala 122:40]
  wire  _T_371 = excMem & memExcept; // @[Mem.scala 123:27]
  wire  _T_372 = _T_370 | _T_371; // @[Mem.scala 122:52]
  wire  _T_373 = _T_372 | excOther; // @[Mem.scala 123:41]
  wire  hasTrap = _T_373 | io_csrHasInt; // @[Mem.scala 123:53]
  wire  _T_375 = ~instIllg; // @[Mem.scala 125:50]
  wire  _T_379 = io_csrMode == 2'h1; // @[Mem.scala 131:33]
  wire [30:0] _T_380 = _T_379 ? 31'h9 : 31'hb; // @[Mem.scala 131:21]
  wire [30:0] _T_381 = _T_353 ? 31'h8 : _T_380; // @[Mem.scala 130:21]
  wire [30:0] _T_382 = memAddr ? 31'h4 : 31'hd; // @[Mem.scala 133:21]
  wire [30:0] _T_383 = memAddr ? 31'h6 : 31'hf; // @[Mem.scala 134:21]
  wire  _T_384 = 4'h9 == io_alu_excType; // @[Mux.scala 68:19]
  wire [30:0] _T_385 = _T_384 ? _T_383 : 31'h0; // @[Mux.scala 68:16]
  wire  _T_386 = 4'h8 == io_alu_excType; // @[Mux.scala 68:19]
  wire [30:0] _T_387 = _T_386 ? _T_382 : _T_385; // @[Mux.scala 68:16]
  wire  _T_388 = 4'h2 == io_alu_excType; // @[Mux.scala 68:19]
  wire [30:0] _T_389 = _T_388 ? 31'h3 : _T_387; // @[Mux.scala 68:16]
  wire  _T_390 = 4'h1 == io_alu_excType; // @[Mux.scala 68:19]
  wire [30:0] cause = _T_390 ? _T_381 : _T_389; // @[Mux.scala 68:16]
  wire [30:0] _T_391 = instAddr ? 31'h0 : cause; // @[Mem.scala 138:22]
  wire [30:0] _T_392 = instIllg ? 31'h2 : _T_391; // @[Mem.scala 137:22]
  wire [31:0] _T_393 = memExcept ? io_alu_reg_data : io_alu_excValue; // @[Mem.scala 143:22]
  wire [31:0] _T_394 = instPage ? io_alu_currentPc : _T_393; // @[Mem.scala 142:22]
  wire  _T_395 = ~stallReq; // @[Mem.scala 147:18]
  wire  _T_396 = flushIc | flushIt; // @[Mem.scala 147:40]
  wire  _T_405 = ~io_csrBusy; // @[Mem.scala 166:26]
  wire  _T_406 = _T_405 & io_alu_valid; // @[Mem.scala 166:38]
  AmoExecute amo ( // @[Mem.scala 55:19]
    .clock(amo_clock),
    .reset(amo_reset),
    .io_op(amo_io_op),
    .io_flush(amo_io_flush),
    .io_ready(amo_io_ready),
    .io_regOpr(amo_io_regOpr),
    .io_regWdata(amo_io_regWdata),
    .io_ramValid(amo_io_ramValid),
    .io_ramWen(amo_io_ramWen),
    .io_ramRdata(amo_io_ramRdata),
    .io_ramWdata(amo_io_ramWdata)
  );
  assign io_stallReq = _T_337 | io_csrBusy; // @[Mem.scala 146:15]
  assign io_flushReq = _T_395 & _T_396; // @[Mem.scala 147:15]
  assign io_flushPc = io_alu_currentPc + 32'h4; // @[Mem.scala 148:15]
  assign io_ram_en = hasTrap ? 1'h0 : en; // @[Mem.scala 151:17]
  assign io_ram_wen = ramWen[3:0]; // @[Mem.scala 152:17]
  assign io_ram_addr = {io_alu_reg_data[31:2],2'h0}; // @[Mem.scala 153:17]
  assign io_ram_wdata = wdata[31:0]; // @[Mem.scala 154:17]
  assign io_flushIc = hasTrap ? 1'h0 : flushIc; // @[Mem.scala 157:15]
  assign io_flushDc = hasTrap ? 1'h0 : flushIc; // @[Mem.scala 158:15]
  assign io_flushIt = hasTrap ? 1'h0 : flushIt; // @[Mem.scala 159:15]
  assign io_flushDt = hasTrap ? 1'h0 : flushIt; // @[Mem.scala 160:15]
  assign io_excMon_addr = {io_alu_reg_data[31:2],2'h0}; // @[Mem.scala 163:19]
  assign io_except_hasTrap = _T_406 & hasTrap; // @[Mem.scala 166:23]
  assign io_except_isSret = _T_352 & _T_375; // @[Mem.scala 167:23]
  assign io_except_isMret = _T_354 & _T_375; // @[Mem.scala 168:23]
  assign io_except_excCause = instPage ? 31'hc : _T_392; // @[Mem.scala 169:23]
  assign io_except_excPc = io_alu_currentPc; // @[Mem.scala 170:23]
  assign io_except_excValue = instIllg ? io_alu_inst : _T_394; // @[Mem.scala 171:23]
  assign io_mem_reg_en = io_alu_reg_en; // @[Mem.scala 174:23]
  assign io_mem_reg_addr = io_alu_reg_addr; // @[Mem.scala 175:23]
  assign io_mem_reg_data = checkExcMon ? {{31'd0}, _T_338} : _T_340; // @[Mem.scala 176:23]
  assign io_mem_reg_load = _T_1 | _T_106; // @[Mem.scala 177:23]
  assign io_mem_memSigned = _T_1 | _T_3; // @[Mem.scala 178:23]
  assign io_mem_memSel = io_alu_reg_data[1:0]; // @[Mem.scala 179:23]
  assign io_mem_memWidth = _T_1 ? 2'h0 : _T_127; // @[Mem.scala 180:23]
  assign io_mem_csr_op = io_alu_csr_op; // @[Mem.scala 181:23]
  assign io_mem_csr_addr = io_alu_csr_addr; // @[Mem.scala 181:23]
  assign io_mem_csr_data = io_alu_csr_data; // @[Mem.scala 181:23]
  assign io_mem_csr_retired = io_alu_csr_retired; // @[Mem.scala 181:23]
  assign io_mem_excMon_addr = {io_alu_reg_data[31:2],2'h0}; // @[Mem.scala 182:23]
  assign io_mem_excMon_set = _T_1 ? 1'h0 : _T_169; // @[Mem.scala 183:23]
  assign io_mem_excMon_clear = _T_331 | _T_332; // @[Mem.scala 184:23]
  assign io_mem_currentPc = io_alu_currentPc; // @[Mem.scala 185:23]
  assign amo_clock = clock;
  assign amo_reset = reset;
  assign amo_io_op = _T_1 ? 4'h0 : _T_211; // @[Mem.scala 56:19]
  assign amo_io_flush = io_flush; // @[Mem.scala 57:19]
  assign amo_io_regOpr = io_alu_lsuData; // @[Mem.scala 58:19]
  assign amo_io_ramValid = io_ram_valid; // @[Mem.scala 59:19]
  assign amo_io_ramRdata = io_ram_rdata; // @[Mem.scala 60:19]
endmodule
module MidStage_3(
  input         clock,
  input         reset,
  input         io_flush,
  input         io_stallPrev,
  input         io_stallNext,
  input         io_prev_reg_en,
  input  [4:0]  io_prev_reg_addr,
  input  [31:0] io_prev_reg_data,
  input         io_prev_reg_load,
  input         io_prev_memSigned,
  input  [1:0]  io_prev_memSel,
  input  [1:0]  io_prev_memWidth,
  input  [2:0]  io_prev_csr_op,
  input  [11:0] io_prev_csr_addr,
  input  [31:0] io_prev_csr_data,
  input         io_prev_csr_retired,
  input  [31:0] io_prev_excMon_addr,
  input         io_prev_excMon_set,
  input         io_prev_excMon_clear,
  input  [31:0] io_prev_currentPc,
  output        io_next_reg_en,
  output [4:0]  io_next_reg_addr,
  output [31:0] io_next_reg_data,
  output        io_next_reg_load,
  output        io_next_memSigned,
  output [1:0]  io_next_memSel,
  output [1:0]  io_next_memWidth,
  output [2:0]  io_next_csr_op,
  output [11:0] io_next_csr_addr,
  output [31:0] io_next_csr_data,
  output        io_next_csr_retired,
  output [31:0] io_next_excMon_addr,
  output        io_next_excMon_set,
  output        io_next_excMon_clear,
  output [31:0] io_next_currentPc
);
  reg  ff_reg_en; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_0;
  reg [4:0] ff_reg_addr; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_1;
  reg [31:0] ff_reg_data; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_2;
  reg  ff_reg_load; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_3;
  reg  ff_memSigned; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_4;
  reg [1:0] ff_memSel; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_5;
  reg [1:0] ff_memWidth; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_6;
  reg [2:0] ff_csr_op; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_7;
  reg [11:0] ff_csr_addr; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_8;
  reg [31:0] ff_csr_data; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_9;
  reg  ff_csr_retired; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_10;
  reg [31:0] ff_excMon_addr; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_11;
  reg  ff_excMon_set; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_12;
  reg  ff_excMon_clear; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_13;
  reg [31:0] ff_currentPc; // @[MidStage.scala 20:19]
  reg [31:0] _RAND_14;
  wire  _T_1 = ~io_stallNext; // @[MidStage.scala 21:38]
  wire  _T_2 = io_stallPrev & _T_1; // @[MidStage.scala 21:35]
  wire  _T_3 = io_flush | _T_2; // @[MidStage.scala 21:18]
  wire  _T_5 = ~io_stallPrev; // @[MidStage.scala 23:15]
  assign io_next_reg_en = ff_reg_en; // @[MidStage.scala 27:11]
  assign io_next_reg_addr = ff_reg_addr; // @[MidStage.scala 27:11]
  assign io_next_reg_data = ff_reg_data; // @[MidStage.scala 27:11]
  assign io_next_reg_load = ff_reg_load; // @[MidStage.scala 27:11]
  assign io_next_memSigned = ff_memSigned; // @[MidStage.scala 27:11]
  assign io_next_memSel = ff_memSel; // @[MidStage.scala 27:11]
  assign io_next_memWidth = ff_memWidth; // @[MidStage.scala 27:11]
  assign io_next_csr_op = ff_csr_op; // @[MidStage.scala 27:11]
  assign io_next_csr_addr = ff_csr_addr; // @[MidStage.scala 27:11]
  assign io_next_csr_data = ff_csr_data; // @[MidStage.scala 27:11]
  assign io_next_csr_retired = ff_csr_retired; // @[MidStage.scala 27:11]
  assign io_next_excMon_addr = ff_excMon_addr; // @[MidStage.scala 27:11]
  assign io_next_excMon_set = ff_excMon_set; // @[MidStage.scala 27:11]
  assign io_next_excMon_clear = ff_excMon_clear; // @[MidStage.scala 27:11]
  assign io_next_currentPc = ff_currentPc; // @[MidStage.scala 27:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  ff_reg_en = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ff_reg_addr = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  ff_reg_data = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  ff_reg_load = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  ff_memSigned = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  ff_memSel = _RAND_5[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  ff_memWidth = _RAND_6[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  ff_csr_op = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  ff_csr_addr = _RAND_8[11:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  ff_csr_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  ff_csr_retired = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  ff_excMon_addr = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  ff_excMon_set = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  ff_excMon_clear = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  ff_currentPc = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      ff_reg_en <= 1'h0;
    end else if (_T_3) begin
      ff_reg_en <= 1'h0;
    end else if (_T_5) begin
      ff_reg_en <= io_prev_reg_en;
    end
    if (reset) begin
      ff_reg_addr <= 5'h0;
    end else if (_T_3) begin
      ff_reg_addr <= 5'h0;
    end else if (_T_5) begin
      ff_reg_addr <= io_prev_reg_addr;
    end
    if (reset) begin
      ff_reg_data <= 32'h0;
    end else if (_T_3) begin
      ff_reg_data <= 32'h0;
    end else if (_T_5) begin
      ff_reg_data <= io_prev_reg_data;
    end
    if (reset) begin
      ff_reg_load <= 1'h0;
    end else if (_T_3) begin
      ff_reg_load <= 1'h0;
    end else if (_T_5) begin
      ff_reg_load <= io_prev_reg_load;
    end
    if (reset) begin
      ff_memSigned <= 1'h0;
    end else if (_T_3) begin
      ff_memSigned <= 1'h0;
    end else if (_T_5) begin
      ff_memSigned <= io_prev_memSigned;
    end
    if (reset) begin
      ff_memSel <= 2'h0;
    end else if (_T_3) begin
      ff_memSel <= 2'h0;
    end else if (_T_5) begin
      ff_memSel <= io_prev_memSel;
    end
    if (reset) begin
      ff_memWidth <= 2'h0;
    end else if (_T_3) begin
      ff_memWidth <= 2'h0;
    end else if (_T_5) begin
      ff_memWidth <= io_prev_memWidth;
    end
    if (reset) begin
      ff_csr_op <= 3'h0;
    end else if (_T_3) begin
      ff_csr_op <= 3'h0;
    end else if (_T_5) begin
      ff_csr_op <= io_prev_csr_op;
    end
    if (reset) begin
      ff_csr_addr <= 12'h0;
    end else if (_T_3) begin
      ff_csr_addr <= 12'h0;
    end else if (_T_5) begin
      ff_csr_addr <= io_prev_csr_addr;
    end
    if (reset) begin
      ff_csr_data <= 32'h0;
    end else if (_T_3) begin
      ff_csr_data <= 32'h0;
    end else if (_T_5) begin
      ff_csr_data <= io_prev_csr_data;
    end
    if (reset) begin
      ff_csr_retired <= 1'h0;
    end else if (_T_3) begin
      ff_csr_retired <= 1'h0;
    end else if (_T_5) begin
      ff_csr_retired <= io_prev_csr_retired;
    end
    if (reset) begin
      ff_excMon_addr <= 32'h0;
    end else if (_T_3) begin
      ff_excMon_addr <= 32'h0;
    end else if (_T_5) begin
      ff_excMon_addr <= io_prev_excMon_addr;
    end
    if (reset) begin
      ff_excMon_set <= 1'h0;
    end else if (_T_3) begin
      ff_excMon_set <= 1'h0;
    end else if (_T_5) begin
      ff_excMon_set <= io_prev_excMon_set;
    end
    if (reset) begin
      ff_excMon_clear <= 1'h0;
    end else if (_T_3) begin
      ff_excMon_clear <= 1'h0;
    end else if (_T_5) begin
      ff_excMon_clear <= io_prev_excMon_clear;
    end
    if (reset) begin
      ff_currentPc <= 32'h0;
    end else if (_T_3) begin
      ff_currentPc <= 32'h0;
    end else if (_T_5) begin
      ff_currentPc <= io_prev_currentPc;
    end
  end
endmodule
module WriteBack(
  input         io_mem_reg_en,
  input  [4:0]  io_mem_reg_addr,
  input  [31:0] io_mem_reg_data,
  input         io_mem_reg_load,
  input         io_mem_memSigned,
  input  [1:0]  io_mem_memSel,
  input  [1:0]  io_mem_memWidth,
  input  [2:0]  io_mem_csr_op,
  input  [11:0] io_mem_csr_addr,
  input  [31:0] io_mem_csr_data,
  input         io_mem_csr_retired,
  input  [31:0] io_mem_excMon_addr,
  input         io_mem_excMon_set,
  input         io_mem_excMon_clear,
  input  [31:0] io_mem_currentPc,
  input  [31:0] io_ramData,
  output        io_reg_en,
  output [4:0]  io_reg_addr,
  output [31:0] io_reg_data,
  output [2:0]  io_csr_op,
  output [11:0] io_csr_addr,
  output [31:0] io_csr_data,
  output        io_csr_retired,
  output [31:0] io_excMon_addr,
  output        io_excMon_set,
  output        io_excMon_clear,
  output        io_debug_regWen,
  output [4:0]  io_debug_regWaddr,
  output [31:0] io_debug_regWdata,
  output [31:0] io_debug_pc
);
  wire [7:0] _T_2 = io_ramData[7:0]; // @[WriteBack.scala 29:15]
  wire [31:0] _T_3 = {{24{_T_2[7]}},_T_2}; // @[WriteBack.scala 30:49]
  wire [31:0] _T_4 = io_mem_memSigned ? _T_3 : {{24'd0}, io_ramData[7:0]}; // @[WriteBack.scala 30:25]
  wire [7:0] _T_7 = io_ramData[15:8]; // @[WriteBack.scala 29:15]
  wire [31:0] _T_8 = {{24{_T_7[7]}},_T_7}; // @[WriteBack.scala 30:49]
  wire [31:0] _T_9 = io_mem_memSigned ? _T_8 : {{24'd0}, io_ramData[15:8]}; // @[WriteBack.scala 30:25]
  wire [7:0] _T_12 = io_ramData[23:16]; // @[WriteBack.scala 29:15]
  wire [31:0] _T_13 = {{24{_T_12[7]}},_T_12}; // @[WriteBack.scala 30:49]
  wire [31:0] _T_14 = io_mem_memSigned ? _T_13 : {{24'd0}, io_ramData[23:16]}; // @[WriteBack.scala 30:25]
  wire [7:0] _T_17 = io_ramData[31:24]; // @[WriteBack.scala 29:15]
  wire [31:0] _T_18 = {{24{_T_17[7]}},_T_17}; // @[WriteBack.scala 30:49]
  wire [31:0] _T_19 = io_mem_memSigned ? _T_18 : {{24'd0}, io_ramData[31:24]}; // @[WriteBack.scala 30:25]
  wire [15:0] _T_22 = io_ramData[15:0]; // @[WriteBack.scala 29:15]
  wire [31:0] _T_23 = {{16{_T_22[15]}},_T_22}; // @[WriteBack.scala 30:49]
  wire [31:0] _T_24 = io_mem_memSigned ? _T_23 : {{16'd0}, io_ramData[15:0]}; // @[WriteBack.scala 30:25]
  wire [15:0] _T_27 = io_ramData[31:16]; // @[WriteBack.scala 29:15]
  wire [31:0] _T_28 = {{16{_T_27[15]}},_T_27}; // @[WriteBack.scala 30:49]
  wire [31:0] _T_29 = io_mem_memSigned ? _T_28 : {{16'd0}, io_ramData[31:16]}; // @[WriteBack.scala 30:25]
  wire [31:0] _T_34 = io_mem_memSigned ? io_ramData : io_ramData; // @[WriteBack.scala 30:25]
  wire  _T_35 = 2'h3 == io_mem_memSel; // @[Mux.scala 68:19]
  wire [31:0] _T_36 = _T_35 ? _T_19 : 32'h0; // @[Mux.scala 68:16]
  wire  _T_37 = 2'h2 == io_mem_memSel; // @[Mux.scala 68:19]
  wire [31:0] _T_38 = _T_37 ? _T_14 : _T_36; // @[Mux.scala 68:16]
  wire  _T_39 = 2'h1 == io_mem_memSel; // @[Mux.scala 68:19]
  wire [31:0] _T_40 = _T_39 ? _T_9 : _T_38; // @[Mux.scala 68:16]
  wire  _T_41 = 2'h0 == io_mem_memSel; // @[Mux.scala 68:19]
  wire [31:0] _T_42 = _T_41 ? _T_4 : _T_40; // @[Mux.scala 68:16]
  wire [31:0] _T_44 = _T_37 ? _T_29 : 32'h0; // @[Mux.scala 68:16]
  wire [31:0] _T_46 = _T_41 ? _T_24 : _T_44; // @[Mux.scala 68:16]
  wire [31:0] _T_48 = _T_41 ? _T_34 : 32'h0; // @[Mux.scala 68:16]
  wire  _T_49 = 2'h2 == io_mem_memWidth; // @[Mux.scala 68:19]
  wire [31:0] _T_50 = _T_49 ? _T_48 : 32'h0; // @[Mux.scala 68:16]
  wire  _T_51 = 2'h1 == io_mem_memWidth; // @[Mux.scala 68:19]
  wire [31:0] _T_52 = _T_51 ? _T_46 : _T_50; // @[Mux.scala 68:16]
  wire  _T_53 = 2'h0 == io_mem_memWidth; // @[Mux.scala 68:19]
  wire [31:0] loadData = _T_53 ? _T_42 : _T_52; // @[Mux.scala 68:16]
  assign io_reg_en = io_mem_reg_en; // @[WriteBack.scala 47:15]
  assign io_reg_addr = io_mem_reg_addr; // @[WriteBack.scala 48:15]
  assign io_reg_data = io_mem_reg_load ? loadData : io_mem_reg_data; // @[WriteBack.scala 49:15]
  assign io_csr_op = io_mem_csr_op; // @[WriteBack.scala 51:15]
  assign io_csr_addr = io_mem_csr_addr; // @[WriteBack.scala 51:15]
  assign io_csr_data = io_mem_csr_data; // @[WriteBack.scala 51:15]
  assign io_csr_retired = io_mem_csr_retired; // @[WriteBack.scala 51:15]
  assign io_excMon_addr = io_mem_excMon_addr; // @[WriteBack.scala 52:15]
  assign io_excMon_set = io_mem_excMon_set; // @[WriteBack.scala 52:15]
  assign io_excMon_clear = io_mem_excMon_clear; // @[WriteBack.scala 52:15]
  assign io_debug_regWen = io_mem_reg_en; // @[WriteBack.scala 55:21]
  assign io_debug_regWaddr = io_mem_reg_addr; // @[WriteBack.scala 56:21]
  assign io_debug_regWdata = io_mem_reg_load ? loadData : io_mem_reg_data; // @[WriteBack.scala 57:21]
  assign io_debug_pc = io_mem_currentPc; // @[WriteBack.scala 58:21]
endmodule
module RegFile(
  input         clock,
  input         reset,
  input         io_read1_en,
  input  [4:0]  io_read1_addr,
  output [31:0] io_read1_data,
  input         io_read2_en,
  input  [4:0]  io_read2_addr,
  output [31:0] io_read2_data,
  input         io_write_en,
  input  [4:0]  io_write_addr,
  input  [31:0] io_write_data
);
  reg [31:0] regfile_0; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_0;
  reg [31:0] regfile_1; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_1;
  reg [31:0] regfile_2; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_2;
  reg [31:0] regfile_3; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_3;
  reg [31:0] regfile_4; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_4;
  reg [31:0] regfile_5; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_5;
  reg [31:0] regfile_6; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_6;
  reg [31:0] regfile_7; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_7;
  reg [31:0] regfile_8; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_8;
  reg [31:0] regfile_9; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_9;
  reg [31:0] regfile_10; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_10;
  reg [31:0] regfile_11; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_11;
  reg [31:0] regfile_12; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_12;
  reg [31:0] regfile_13; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_13;
  reg [31:0] regfile_14; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_14;
  reg [31:0] regfile_15; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_15;
  reg [31:0] regfile_16; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_16;
  reg [31:0] regfile_17; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_17;
  reg [31:0] regfile_18; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_18;
  reg [31:0] regfile_19; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_19;
  reg [31:0] regfile_20; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_20;
  reg [31:0] regfile_21; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_21;
  reg [31:0] regfile_22; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_22;
  reg [31:0] regfile_23; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_23;
  reg [31:0] regfile_24; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_24;
  reg [31:0] regfile_25; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_25;
  reg [31:0] regfile_26; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_26;
  reg [31:0] regfile_27; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_27;
  reg [31:0] regfile_28; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_28;
  reg [31:0] regfile_29; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_29;
  reg [31:0] regfile_30; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_30;
  reg [31:0] regfile_31; // @[RegFile.scala 17:24]
  reg [31:0] _RAND_31;
  wire [31:0] _GEN_1 = 5'h1 == io_read1_addr ? regfile_1 : regfile_0; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_2 = 5'h2 == io_read1_addr ? regfile_2 : _GEN_1; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_3 = 5'h3 == io_read1_addr ? regfile_3 : _GEN_2; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_4 = 5'h4 == io_read1_addr ? regfile_4 : _GEN_3; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_5 = 5'h5 == io_read1_addr ? regfile_5 : _GEN_4; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_6 = 5'h6 == io_read1_addr ? regfile_6 : _GEN_5; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_7 = 5'h7 == io_read1_addr ? regfile_7 : _GEN_6; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_8 = 5'h8 == io_read1_addr ? regfile_8 : _GEN_7; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_9 = 5'h9 == io_read1_addr ? regfile_9 : _GEN_8; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_10 = 5'ha == io_read1_addr ? regfile_10 : _GEN_9; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_11 = 5'hb == io_read1_addr ? regfile_11 : _GEN_10; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_12 = 5'hc == io_read1_addr ? regfile_12 : _GEN_11; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_13 = 5'hd == io_read1_addr ? regfile_13 : _GEN_12; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_14 = 5'he == io_read1_addr ? regfile_14 : _GEN_13; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_15 = 5'hf == io_read1_addr ? regfile_15 : _GEN_14; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_16 = 5'h10 == io_read1_addr ? regfile_16 : _GEN_15; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_17 = 5'h11 == io_read1_addr ? regfile_17 : _GEN_16; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_18 = 5'h12 == io_read1_addr ? regfile_18 : _GEN_17; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_19 = 5'h13 == io_read1_addr ? regfile_19 : _GEN_18; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_20 = 5'h14 == io_read1_addr ? regfile_20 : _GEN_19; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_21 = 5'h15 == io_read1_addr ? regfile_21 : _GEN_20; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_22 = 5'h16 == io_read1_addr ? regfile_22 : _GEN_21; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_23 = 5'h17 == io_read1_addr ? regfile_23 : _GEN_22; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_24 = 5'h18 == io_read1_addr ? regfile_24 : _GEN_23; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_25 = 5'h19 == io_read1_addr ? regfile_25 : _GEN_24; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_26 = 5'h1a == io_read1_addr ? regfile_26 : _GEN_25; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_27 = 5'h1b == io_read1_addr ? regfile_27 : _GEN_26; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_28 = 5'h1c == io_read1_addr ? regfile_28 : _GEN_27; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_29 = 5'h1d == io_read1_addr ? regfile_29 : _GEN_28; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_30 = 5'h1e == io_read1_addr ? regfile_30 : _GEN_29; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_31 = 5'h1f == io_read1_addr ? regfile_31 : _GEN_30; // @[RegFile.scala 20:23]
  wire [31:0] _GEN_33 = 5'h1 == io_read2_addr ? regfile_1 : regfile_0; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_34 = 5'h2 == io_read2_addr ? regfile_2 : _GEN_33; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_35 = 5'h3 == io_read2_addr ? regfile_3 : _GEN_34; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_36 = 5'h4 == io_read2_addr ? regfile_4 : _GEN_35; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_37 = 5'h5 == io_read2_addr ? regfile_5 : _GEN_36; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_38 = 5'h6 == io_read2_addr ? regfile_6 : _GEN_37; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_39 = 5'h7 == io_read2_addr ? regfile_7 : _GEN_38; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_40 = 5'h8 == io_read2_addr ? regfile_8 : _GEN_39; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_41 = 5'h9 == io_read2_addr ? regfile_9 : _GEN_40; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_42 = 5'ha == io_read2_addr ? regfile_10 : _GEN_41; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_43 = 5'hb == io_read2_addr ? regfile_11 : _GEN_42; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_44 = 5'hc == io_read2_addr ? regfile_12 : _GEN_43; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_45 = 5'hd == io_read2_addr ? regfile_13 : _GEN_44; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_46 = 5'he == io_read2_addr ? regfile_14 : _GEN_45; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_47 = 5'hf == io_read2_addr ? regfile_15 : _GEN_46; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_48 = 5'h10 == io_read2_addr ? regfile_16 : _GEN_47; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_49 = 5'h11 == io_read2_addr ? regfile_17 : _GEN_48; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_50 = 5'h12 == io_read2_addr ? regfile_18 : _GEN_49; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_51 = 5'h13 == io_read2_addr ? regfile_19 : _GEN_50; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_52 = 5'h14 == io_read2_addr ? regfile_20 : _GEN_51; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_53 = 5'h15 == io_read2_addr ? regfile_21 : _GEN_52; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_54 = 5'h16 == io_read2_addr ? regfile_22 : _GEN_53; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_55 = 5'h17 == io_read2_addr ? regfile_23 : _GEN_54; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_56 = 5'h18 == io_read2_addr ? regfile_24 : _GEN_55; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_57 = 5'h19 == io_read2_addr ? regfile_25 : _GEN_56; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_58 = 5'h1a == io_read2_addr ? regfile_26 : _GEN_57; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_59 = 5'h1b == io_read2_addr ? regfile_27 : _GEN_58; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_60 = 5'h1c == io_read2_addr ? regfile_28 : _GEN_59; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_61 = 5'h1d == io_read2_addr ? regfile_29 : _GEN_60; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_62 = 5'h1e == io_read2_addr ? regfile_30 : _GEN_61; // @[RegFile.scala 21:23]
  wire [31:0] _GEN_63 = 5'h1f == io_read2_addr ? regfile_31 : _GEN_62; // @[RegFile.scala 21:23]
  wire  _T_3 = io_write_addr != 5'h0; // @[RegFile.scala 24:38]
  wire  _T_4 = io_write_en & _T_3; // @[RegFile.scala 24:21]
  assign io_read1_data = io_read1_en ? _GEN_31 : 32'h0; // @[RegFile.scala 20:17]
  assign io_read2_data = io_read2_en ? _GEN_63 : 32'h0; // @[RegFile.scala 21:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regfile_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  regfile_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  regfile_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  regfile_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  regfile_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  regfile_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  regfile_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  regfile_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  regfile_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  regfile_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  regfile_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  regfile_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  regfile_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  regfile_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  regfile_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  regfile_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  regfile_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  regfile_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  regfile_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  regfile_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  regfile_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  regfile_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  regfile_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  regfile_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  regfile_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  regfile_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  regfile_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  regfile_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  regfile_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  regfile_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  regfile_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  regfile_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      regfile_0 <= 32'h0;
    end else if (_T_4) begin
      if (5'h0 == io_write_addr) begin
        regfile_0 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_1 <= 32'h0;
    end else if (_T_4) begin
      if (5'h1 == io_write_addr) begin
        regfile_1 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_2 <= 32'h0;
    end else if (_T_4) begin
      if (5'h2 == io_write_addr) begin
        regfile_2 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_3 <= 32'h0;
    end else if (_T_4) begin
      if (5'h3 == io_write_addr) begin
        regfile_3 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_4 <= 32'h0;
    end else if (_T_4) begin
      if (5'h4 == io_write_addr) begin
        regfile_4 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_5 <= 32'h0;
    end else if (_T_4) begin
      if (5'h5 == io_write_addr) begin
        regfile_5 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_6 <= 32'h0;
    end else if (_T_4) begin
      if (5'h6 == io_write_addr) begin
        regfile_6 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_7 <= 32'h0;
    end else if (_T_4) begin
      if (5'h7 == io_write_addr) begin
        regfile_7 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_8 <= 32'h0;
    end else if (_T_4) begin
      if (5'h8 == io_write_addr) begin
        regfile_8 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_9 <= 32'h0;
    end else if (_T_4) begin
      if (5'h9 == io_write_addr) begin
        regfile_9 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_10 <= 32'h0;
    end else if (_T_4) begin
      if (5'ha == io_write_addr) begin
        regfile_10 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_11 <= 32'h0;
    end else if (_T_4) begin
      if (5'hb == io_write_addr) begin
        regfile_11 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_12 <= 32'h0;
    end else if (_T_4) begin
      if (5'hc == io_write_addr) begin
        regfile_12 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_13 <= 32'h0;
    end else if (_T_4) begin
      if (5'hd == io_write_addr) begin
        regfile_13 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_14 <= 32'h0;
    end else if (_T_4) begin
      if (5'he == io_write_addr) begin
        regfile_14 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_15 <= 32'h0;
    end else if (_T_4) begin
      if (5'hf == io_write_addr) begin
        regfile_15 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_16 <= 32'h0;
    end else if (_T_4) begin
      if (5'h10 == io_write_addr) begin
        regfile_16 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_17 <= 32'h0;
    end else if (_T_4) begin
      if (5'h11 == io_write_addr) begin
        regfile_17 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_18 <= 32'h0;
    end else if (_T_4) begin
      if (5'h12 == io_write_addr) begin
        regfile_18 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_19 <= 32'h0;
    end else if (_T_4) begin
      if (5'h13 == io_write_addr) begin
        regfile_19 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_20 <= 32'h0;
    end else if (_T_4) begin
      if (5'h14 == io_write_addr) begin
        regfile_20 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_21 <= 32'h0;
    end else if (_T_4) begin
      if (5'h15 == io_write_addr) begin
        regfile_21 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_22 <= 32'h0;
    end else if (_T_4) begin
      if (5'h16 == io_write_addr) begin
        regfile_22 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_23 <= 32'h0;
    end else if (_T_4) begin
      if (5'h17 == io_write_addr) begin
        regfile_23 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_24 <= 32'h0;
    end else if (_T_4) begin
      if (5'h18 == io_write_addr) begin
        regfile_24 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_25 <= 32'h0;
    end else if (_T_4) begin
      if (5'h19 == io_write_addr) begin
        regfile_25 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_26 <= 32'h0;
    end else if (_T_4) begin
      if (5'h1a == io_write_addr) begin
        regfile_26 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_27 <= 32'h0;
    end else if (_T_4) begin
      if (5'h1b == io_write_addr) begin
        regfile_27 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_28 <= 32'h0;
    end else if (_T_4) begin
      if (5'h1c == io_write_addr) begin
        regfile_28 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_29 <= 32'h0;
    end else if (_T_4) begin
      if (5'h1d == io_write_addr) begin
        regfile_29 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_30 <= 32'h0;
    end else if (_T_4) begin
      if (5'h1e == io_write_addr) begin
        regfile_30 <= io_write_data;
      end
    end
    if (reset) begin
      regfile_31 <= 32'h0;
    end else if (_T_4) begin
      if (5'h1f == io_write_addr) begin
        regfile_31 <= io_write_data;
      end
    end
  end
endmodule
module CsrFile(
  input         clock,
  input         reset,
  input  [2:0]  io_read_op,
  output        io_read_valid,
  input  [11:0] io_read_addr,
  output [31:0] io_read_data,
  input  [2:0]  io_write_op,
  input  [11:0] io_write_addr,
  input  [31:0] io_write_data,
  input         io_write_retired,
  input         io_irq_timer,
  input         io_irq_soft,
  input         io_irq_extern,
  input         io_except_hasTrap,
  input         io_except_isSret,
  input         io_except_isMret,
  input  [30:0] io_except_excCause,
  input  [31:0] io_except_excPc,
  input  [31:0] io_except_excValue,
  output        io_hasInt,
  output        io_busy,
  output [1:0]  io_mode,
  output [31:0] io_sepc,
  output [31:0] io_mepc,
  output [31:0] io_trapVec,
  output        io_pageEn,
  output [21:0] io_basePpn,
  output        io_sum
);
  reg [1:0] mode; // @[CsrFile.scala 39:26]
  reg [31:0] _RAND_0;
  reg  mstatus_sum; // @[CsrFile.scala 42:26]
  reg [31:0] _RAND_1;
  reg [1:0] mstatus_mpp; // @[CsrFile.scala 42:26]
  reg [31:0] _RAND_2;
  reg  mstatus_spp; // @[CsrFile.scala 42:26]
  reg [31:0] _RAND_3;
  reg  mstatus_mpie; // @[CsrFile.scala 42:26]
  reg [31:0] _RAND_4;
  reg  mstatus_spie; // @[CsrFile.scala 42:26]
  reg [31:0] _RAND_5;
  reg  mstatus_mie; // @[CsrFile.scala 42:26]
  reg [31:0] _RAND_6;
  reg  mstatus_sie; // @[CsrFile.scala 42:26]
  reg [31:0] _RAND_7;
  reg [31:0] medeleg_data; // @[CsrFile.scala 44:26]
  reg [31:0] _RAND_8;
  reg [31:0] mideleg_data; // @[CsrFile.scala 45:26]
  reg [31:0] _RAND_9;
  reg  mie_meie; // @[CsrFile.scala 46:26]
  reg [31:0] _RAND_10;
  reg  mie_seie; // @[CsrFile.scala 46:26]
  reg [31:0] _RAND_11;
  reg  mie_mtie; // @[CsrFile.scala 46:26]
  reg [31:0] _RAND_12;
  reg  mie_stie; // @[CsrFile.scala 46:26]
  reg [31:0] _RAND_13;
  reg  mie_msie; // @[CsrFile.scala 46:26]
  reg [31:0] _RAND_14;
  reg  mie_ssie; // @[CsrFile.scala 46:26]
  reg [31:0] _RAND_15;
  reg [29:0] mtvec_base; // @[CsrFile.scala 47:26]
  reg [31:0] _RAND_16;
  reg [1:0] mtvec_mode; // @[CsrFile.scala 47:26]
  reg [31:0] _RAND_17;
  reg [31:0] mscratch_data; // @[CsrFile.scala 48:26]
  reg [31:0] _RAND_18;
  reg [31:0] mepc_data; // @[CsrFile.scala 49:26]
  reg [31:0] _RAND_19;
  reg  mcause_int; // @[CsrFile.scala 50:26]
  reg [31:0] _RAND_20;
  reg [30:0] mcause_code; // @[CsrFile.scala 50:26]
  reg [31:0] _RAND_21;
  reg [31:0] mtval_data; // @[CsrFile.scala 51:26]
  reg [31:0] _RAND_22;
  reg  mipReal_seip; // @[CsrFile.scala 52:26]
  reg [31:0] _RAND_23;
  reg  mipReal_stip; // @[CsrFile.scala 52:26]
  reg [31:0] _RAND_24;
  reg  mipReal_ssip; // @[CsrFile.scala 52:26]
  reg [31:0] _RAND_25;
  reg [63:0] mcycle_data; // @[CsrFile.scala 54:26]
  reg [63:0] _RAND_26;
  reg [63:0] minstret_data; // @[CsrFile.scala 55:26]
  reg [63:0] _RAND_27;
  wire [10:0] _T_20 = {2'h0,mstatus_spp,mstatus_mpie,1'h0,mstatus_spie,1'h0,mstatus_mie,1'h0,mstatus_sie,1'h0}; // @[CSR.scala 31:18]
  wire [31:0] _T_31 = {13'h0,mstatus_sum,1'h0,2'h0,2'h0,mstatus_mpp,_T_20}; // @[CSR.scala 31:18]
  wire  sstatus_sum = _T_31[18]; // @[CSR.scala 56:18]
  wire  sstatus_spp = _T_31[8]; // @[CSR.scala 57:18]
  wire  sstatus_spie = _T_31[5]; // @[CSR.scala 58:18]
  wire  sstatus_sie = _T_31[1]; // @[CSR.scala 59:18]
  wire [5:0] _T_40 = {mie_stie,1'h0,mie_msie,1'h0,mie_ssie,1'h0}; // @[CSR.scala 31:18]
  wire [31:0] _T_47 = {20'h0,mie_meie,1'h0,mie_seie,1'h0,mie_mtie,1'h0,_T_40}; // @[CSR.scala 31:18]
  wire  sie_seie = _T_47[9]; // @[CSR.scala 81:18]
  wire  sie_stie = _T_47[5]; // @[CSR.scala 82:18]
  wire  sie_ssie = _T_47[1]; // @[CSR.scala 83:18]
  reg [29:0] stvec_base; // @[CsrFile.scala 59:26]
  reg [31:0] _RAND_28;
  reg [1:0] stvec_mode; // @[CsrFile.scala 59:26]
  reg [31:0] _RAND_29;
  reg [31:0] sscratch_data; // @[CsrFile.scala 60:26]
  reg [31:0] _RAND_30;
  reg [31:0] sepc_data; // @[CsrFile.scala 61:26]
  reg [31:0] _RAND_31;
  reg  scause_int; // @[CsrFile.scala 62:26]
  reg [31:0] _RAND_32;
  reg [30:0] scause_code; // @[CsrFile.scala 62:26]
  reg [31:0] _RAND_33;
  reg [31:0] stval_data; // @[CsrFile.scala 63:26]
  reg [31:0] _RAND_34;
  reg  satp_mode; // @[CsrFile.scala 64:26]
  reg [31:0] _RAND_35;
  reg [21:0] satp_ppn; // @[CsrFile.scala 64:26]
  reg [31:0] _RAND_36;
  wire [8:0] _T_66 = {sstatus_spp,2'h0,sstatus_spie,1'h0,2'h0,sstatus_sie,1'h0}; // @[CsrFile.scala 79:48]
  wire [31:0] _T_74 = {12'h0,1'h0,sstatus_sum,9'h0,_T_66}; // @[CsrFile.scala 79:48]
  wire [31:0] _T_82 = {22'h0,sie_seie,1'h0,2'h0,sie_stie,3'h0,sie_ssie,1'h0}; // @[CsrFile.scala 80:44]
  wire [31:0] _T_83 = {stvec_base,stvec_mode}; // @[CsrFile.scala 81:46]
  wire [31:0] _T_84 = {scause_int,scause_code}; // @[CsrFile.scala 85:47]
  wire  mip_ssip = mipReal_ssip | io_irq_soft; // @[CsrFile.scala 191:28]
  wire  mip_stip = mipReal_stip | io_irq_timer; // @[CsrFile.scala 189:28]
  wire  mip_seip = mipReal_seip | io_irq_extern; // @[CsrFile.scala 187:28]
  wire [31:0] _T_92 = {22'h0,mip_seip,1'h0,2'h0,mip_stip,3'h0,mip_ssip,1'h0}; // @[CsrFile.scala 87:44]
  wire [31:0] _T_94 = {satp_mode,9'h0,satp_ppn}; // @[CsrFile.scala 88:45]
  wire [31:0] _T_129 = {mtvec_base,mtvec_mode}; // @[CsrFile.scala 98:46]
  wire [31:0] _T_130 = {mcause_int,mcause_code}; // @[CsrFile.scala 102:47]
  wire [5:0] _T_135 = {mip_stip,1'h0,io_irq_soft,1'h0,mip_ssip,1'h0}; // @[CsrFile.scala 104:44]
  wire [31:0] _T_142 = {20'h0,io_irq_extern,1'h0,mip_seip,1'h0,io_irq_timer,1'h0,_T_135}; // @[CsrFile.scala 104:44]
  wire  _T_148 = 12'hc00 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_150 = 12'hc02 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_152 = 12'hc80 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_154 = 12'hc82 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_156 = 12'h100 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_158 = 12'h104 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_160 = 12'h105 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_162 = 12'h106 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_164 = 12'h140 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_166 = 12'h141 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_168 = 12'h142 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_170 = 12'h143 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_172 = 12'h144 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_174 = 12'h180 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_176 = 12'hf11 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_178 = 12'hf12 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_180 = 12'hf13 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_182 = 12'hf14 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_184 = 12'h300 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_186 = 12'h301 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_188 = 12'h302 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_190 = 12'h303 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_192 = 12'h304 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_194 = 12'h305 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_196 = 12'h306 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_198 = 12'h340 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_200 = 12'h341 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_202 = 12'h342 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_204 = 12'h343 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_206 = 12'h344 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_208 = 12'h3a0 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_210 = 12'h3a1 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_212 = 12'h3a2 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_214 = 12'h3a3 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_216 = 12'h3b0 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_218 = 12'h3b1 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_220 = 12'h3b2 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_222 = 12'h3b3 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_224 = 12'h3b4 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_226 = 12'h3b5 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_228 = 12'h3b6 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_230 = 12'h3b7 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_232 = 12'h3b8 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_234 = 12'h3b9 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_236 = 12'h3ba == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_238 = 12'h3bb == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_240 = 12'h3bc == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_242 = 12'h3bd == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_244 = 12'h3be == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_246 = 12'h3bf == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_248 = 12'hb00 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_250 = 12'hb02 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_252 = 12'hb80 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_254 = 12'hb82 == io_read_addr; // @[Lookup.scala 31:38]
  wire  _T_256 = 12'h320 == io_read_addr; // @[Lookup.scala 31:38]
  wire [31:0] _T_258 = _T_254 ? minstret_data[63:32] : 32'h0; // @[Lookup.scala 33:37]
  wire [31:0] _T_259 = _T_252 ? mcycle_data[63:32] : _T_258; // @[Lookup.scala 33:37]
  wire [31:0] _T_260 = _T_250 ? minstret_data[31:0] : _T_259; // @[Lookup.scala 33:37]
  wire [31:0] _T_261 = _T_248 ? mcycle_data[31:0] : _T_260; // @[Lookup.scala 33:37]
  wire [31:0] _T_262 = _T_246 ? 32'h0 : _T_261; // @[Lookup.scala 33:37]
  wire [31:0] _T_263 = _T_244 ? 32'h0 : _T_262; // @[Lookup.scala 33:37]
  wire [31:0] _T_264 = _T_242 ? 32'h0 : _T_263; // @[Lookup.scala 33:37]
  wire [31:0] _T_265 = _T_240 ? 32'h0 : _T_264; // @[Lookup.scala 33:37]
  wire [31:0] _T_266 = _T_238 ? 32'h0 : _T_265; // @[Lookup.scala 33:37]
  wire [31:0] _T_267 = _T_236 ? 32'h0 : _T_266; // @[Lookup.scala 33:37]
  wire [31:0] _T_268 = _T_234 ? 32'h0 : _T_267; // @[Lookup.scala 33:37]
  wire [31:0] _T_269 = _T_232 ? 32'h0 : _T_268; // @[Lookup.scala 33:37]
  wire [31:0] _T_270 = _T_230 ? 32'h0 : _T_269; // @[Lookup.scala 33:37]
  wire [31:0] _T_271 = _T_228 ? 32'h0 : _T_270; // @[Lookup.scala 33:37]
  wire [31:0] _T_272 = _T_226 ? 32'h0 : _T_271; // @[Lookup.scala 33:37]
  wire [31:0] _T_273 = _T_224 ? 32'h0 : _T_272; // @[Lookup.scala 33:37]
  wire [31:0] _T_274 = _T_222 ? 32'h0 : _T_273; // @[Lookup.scala 33:37]
  wire [31:0] _T_275 = _T_220 ? 32'h0 : _T_274; // @[Lookup.scala 33:37]
  wire [31:0] _T_276 = _T_218 ? 32'h0 : _T_275; // @[Lookup.scala 33:37]
  wire [31:0] _T_277 = _T_216 ? 32'h0 : _T_276; // @[Lookup.scala 33:37]
  wire [31:0] _T_278 = _T_214 ? 32'h0 : _T_277; // @[Lookup.scala 33:37]
  wire [31:0] _T_279 = _T_212 ? 32'h0 : _T_278; // @[Lookup.scala 33:37]
  wire [31:0] _T_280 = _T_210 ? 32'h0 : _T_279; // @[Lookup.scala 33:37]
  wire [31:0] _T_281 = _T_208 ? 32'h0 : _T_280; // @[Lookup.scala 33:37]
  wire [31:0] _T_282 = _T_206 ? _T_142 : _T_281; // @[Lookup.scala 33:37]
  wire [31:0] _T_283 = _T_204 ? mtval_data : _T_282; // @[Lookup.scala 33:37]
  wire [31:0] _T_284 = _T_202 ? _T_130 : _T_283; // @[Lookup.scala 33:37]
  wire [31:0] _T_285 = _T_200 ? mepc_data : _T_284; // @[Lookup.scala 33:37]
  wire [31:0] _T_286 = _T_198 ? mscratch_data : _T_285; // @[Lookup.scala 33:37]
  wire [31:0] _T_287 = _T_196 ? 32'h0 : _T_286; // @[Lookup.scala 33:37]
  wire [31:0] _T_288 = _T_194 ? _T_129 : _T_287; // @[Lookup.scala 33:37]
  wire [31:0] _T_289 = _T_192 ? _T_47 : _T_288; // @[Lookup.scala 33:37]
  wire [31:0] _T_290 = _T_190 ? mideleg_data : _T_289; // @[Lookup.scala 33:37]
  wire [31:0] _T_291 = _T_188 ? medeleg_data : _T_290; // @[Lookup.scala 33:37]
  wire [31:0] _T_292 = _T_186 ? 32'h40141101 : _T_291; // @[Lookup.scala 33:37]
  wire [31:0] _T_293 = _T_184 ? _T_31 : _T_292; // @[Lookup.scala 33:37]
  wire [31:0] _T_294 = _T_182 ? 32'h0 : _T_293; // @[Lookup.scala 33:37]
  wire [31:0] _T_295 = _T_180 ? 32'h0 : _T_294; // @[Lookup.scala 33:37]
  wire [31:0] _T_296 = _T_178 ? 32'h0 : _T_295; // @[Lookup.scala 33:37]
  wire [31:0] _T_297 = _T_176 ? 32'h0 : _T_296; // @[Lookup.scala 33:37]
  wire [31:0] _T_298 = _T_174 ? _T_94 : _T_297; // @[Lookup.scala 33:37]
  wire [31:0] _T_299 = _T_172 ? _T_92 : _T_298; // @[Lookup.scala 33:37]
  wire [31:0] _T_300 = _T_170 ? stval_data : _T_299; // @[Lookup.scala 33:37]
  wire [31:0] _T_301 = _T_168 ? _T_84 : _T_300; // @[Lookup.scala 33:37]
  wire [31:0] _T_302 = _T_166 ? sepc_data : _T_301; // @[Lookup.scala 33:37]
  wire [31:0] _T_303 = _T_164 ? sscratch_data : _T_302; // @[Lookup.scala 33:37]
  wire [31:0] _T_304 = _T_162 ? 32'h0 : _T_303; // @[Lookup.scala 33:37]
  wire [31:0] _T_305 = _T_160 ? _T_83 : _T_304; // @[Lookup.scala 33:37]
  wire [31:0] _T_306 = _T_158 ? _T_82 : _T_305; // @[Lookup.scala 33:37]
  wire [31:0] _T_307 = _T_156 ? _T_74 : _T_306; // @[Lookup.scala 33:37]
  wire [31:0] _T_308 = _T_154 ? minstret_data[63:32] : _T_307; // @[Lookup.scala 33:37]
  wire [31:0] _T_309 = _T_152 ? mcycle_data[63:32] : _T_308; // @[Lookup.scala 33:37]
  wire [31:0] _T_310 = _T_150 ? minstret_data[31:0] : _T_309; // @[Lookup.scala 33:37]
  wire  _T_312 = _T_254 | _T_256; // @[Lookup.scala 33:37]
  wire  _T_313 = _T_252 | _T_312; // @[Lookup.scala 33:37]
  wire  _T_314 = _T_250 | _T_313; // @[Lookup.scala 33:37]
  wire  _T_315 = _T_248 | _T_314; // @[Lookup.scala 33:37]
  wire  _T_316 = _T_246 | _T_315; // @[Lookup.scala 33:37]
  wire  _T_317 = _T_244 | _T_316; // @[Lookup.scala 33:37]
  wire  _T_318 = _T_242 | _T_317; // @[Lookup.scala 33:37]
  wire  _T_319 = _T_240 | _T_318; // @[Lookup.scala 33:37]
  wire  _T_320 = _T_238 | _T_319; // @[Lookup.scala 33:37]
  wire  _T_321 = _T_236 | _T_320; // @[Lookup.scala 33:37]
  wire  _T_322 = _T_234 | _T_321; // @[Lookup.scala 33:37]
  wire  _T_323 = _T_232 | _T_322; // @[Lookup.scala 33:37]
  wire  _T_324 = _T_230 | _T_323; // @[Lookup.scala 33:37]
  wire  _T_325 = _T_228 | _T_324; // @[Lookup.scala 33:37]
  wire  _T_326 = _T_226 | _T_325; // @[Lookup.scala 33:37]
  wire  _T_327 = _T_224 | _T_326; // @[Lookup.scala 33:37]
  wire  _T_328 = _T_222 | _T_327; // @[Lookup.scala 33:37]
  wire  _T_329 = _T_220 | _T_328; // @[Lookup.scala 33:37]
  wire  _T_330 = _T_218 | _T_329; // @[Lookup.scala 33:37]
  wire  _T_331 = _T_216 | _T_330; // @[Lookup.scala 33:37]
  wire  _T_332 = _T_214 | _T_331; // @[Lookup.scala 33:37]
  wire  _T_333 = _T_212 | _T_332; // @[Lookup.scala 33:37]
  wire  _T_334 = _T_210 | _T_333; // @[Lookup.scala 33:37]
  wire  _T_335 = _T_208 | _T_334; // @[Lookup.scala 33:37]
  wire  _T_336 = _T_206 | _T_335; // @[Lookup.scala 33:37]
  wire  _T_337 = _T_204 | _T_336; // @[Lookup.scala 33:37]
  wire  _T_338 = _T_202 | _T_337; // @[Lookup.scala 33:37]
  wire  _T_339 = _T_200 | _T_338; // @[Lookup.scala 33:37]
  wire  _T_340 = _T_198 | _T_339; // @[Lookup.scala 33:37]
  wire  _T_341 = _T_196 | _T_340; // @[Lookup.scala 33:37]
  wire  _T_342 = _T_194 | _T_341; // @[Lookup.scala 33:37]
  wire  _T_343 = _T_192 | _T_342; // @[Lookup.scala 33:37]
  wire  _T_344 = _T_190 | _T_343; // @[Lookup.scala 33:37]
  wire  _T_345 = _T_188 | _T_344; // @[Lookup.scala 33:37]
  wire  _T_346 = _T_186 | _T_345; // @[Lookup.scala 33:37]
  wire  _T_347 = _T_184 | _T_346; // @[Lookup.scala 33:37]
  wire  _T_348 = _T_182 | _T_347; // @[Lookup.scala 33:37]
  wire  _T_349 = _T_180 | _T_348; // @[Lookup.scala 33:37]
  wire  _T_350 = _T_178 | _T_349; // @[Lookup.scala 33:37]
  wire  _T_351 = _T_176 | _T_350; // @[Lookup.scala 33:37]
  wire  _T_352 = _T_174 | _T_351; // @[Lookup.scala 33:37]
  wire  _T_353 = _T_172 | _T_352; // @[Lookup.scala 33:37]
  wire  _T_354 = _T_170 | _T_353; // @[Lookup.scala 33:37]
  wire  _T_355 = _T_168 | _T_354; // @[Lookup.scala 33:37]
  wire  _T_356 = _T_166 | _T_355; // @[Lookup.scala 33:37]
  wire  _T_357 = _T_164 | _T_356; // @[Lookup.scala 33:37]
  wire  _T_358 = _T_162 | _T_357; // @[Lookup.scala 33:37]
  wire  _T_359 = _T_160 | _T_358; // @[Lookup.scala 33:37]
  wire  _T_360 = _T_158 | _T_359; // @[Lookup.scala 33:37]
  wire  _T_361 = _T_156 | _T_360; // @[Lookup.scala 33:37]
  wire  _T_362 = _T_154 | _T_361; // @[Lookup.scala 33:37]
  wire  _T_363 = _T_152 | _T_362; // @[Lookup.scala 33:37]
  wire  _T_364 = _T_150 | _T_363; // @[Lookup.scala 33:37]
  wire  readable = _T_148 | _T_364; // @[Lookup.scala 33:37]
  wire  _T_402 = _T_182 ? 1'h0 : _T_347; // @[Lookup.scala 33:37]
  wire  _T_403 = _T_180 ? 1'h0 : _T_402; // @[Lookup.scala 33:37]
  wire  _T_404 = _T_178 ? 1'h0 : _T_403; // @[Lookup.scala 33:37]
  wire  _T_405 = _T_176 ? 1'h0 : _T_404; // @[Lookup.scala 33:37]
  wire  _T_406 = _T_174 | _T_405; // @[Lookup.scala 33:37]
  wire  _T_407 = _T_172 | _T_406; // @[Lookup.scala 33:37]
  wire  _T_408 = _T_170 | _T_407; // @[Lookup.scala 33:37]
  wire  _T_409 = _T_168 | _T_408; // @[Lookup.scala 33:37]
  wire  _T_410 = _T_166 | _T_409; // @[Lookup.scala 33:37]
  wire  _T_411 = _T_164 | _T_410; // @[Lookup.scala 33:37]
  wire  _T_412 = _T_162 | _T_411; // @[Lookup.scala 33:37]
  wire  _T_413 = _T_160 | _T_412; // @[Lookup.scala 33:37]
  wire  _T_414 = _T_158 | _T_413; // @[Lookup.scala 33:37]
  wire  _T_415 = _T_156 | _T_414; // @[Lookup.scala 33:37]
  wire  _T_416 = _T_154 ? 1'h0 : _T_415; // @[Lookup.scala 33:37]
  wire  _T_417 = _T_152 ? 1'h0 : _T_416; // @[Lookup.scala 33:37]
  wire  _T_418 = _T_150 ? 1'h0 : _T_417; // @[Lookup.scala 33:37]
  wire  writable = _T_148 ? 1'h0 : _T_418; // @[Lookup.scala 33:37]
  wire  _T_419 = readable & writable; // @[CsrFile.scala 138:26]
  wire  _T_422 = 3'h5 == io_read_op; // @[Mux.scala 68:19]
  wire  _T_423 = _T_422 & _T_419; // @[Mux.scala 68:16]
  wire  _T_424 = 3'h4 == io_read_op; // @[Mux.scala 68:19]
  wire  _T_425 = _T_424 ? _T_419 : _T_423; // @[Mux.scala 68:16]
  wire  _T_426 = 3'h3 == io_read_op; // @[Mux.scala 68:19]
  wire  _T_427 = _T_426 ? _T_419 : _T_425; // @[Mux.scala 68:16]
  wire  _T_428 = 3'h2 == io_read_op; // @[Mux.scala 68:19]
  wire  _T_429 = _T_428 ? writable : _T_427; // @[Mux.scala 68:16]
  wire  _T_430 = 3'h1 == io_read_op; // @[Mux.scala 68:19]
  wire  readValid = _T_430 ? readable : _T_429; // @[Mux.scala 68:16]
  wire  modeValid = io_read_addr[9:8] <= mode; // @[CsrFile.scala 142:38]
  wire  _T_433 = 12'hc00 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_435 = 12'hc02 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_437 = 12'hc80 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_439 = 12'hc82 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_441 = 12'h100 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_443 = 12'h104 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_445 = 12'h105 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_447 = 12'h106 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_449 = 12'h140 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_451 = 12'h141 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_453 = 12'h142 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_455 = 12'h143 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_457 = 12'h144 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_459 = 12'h180 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_461 = 12'hf11 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_463 = 12'hf12 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_465 = 12'hf13 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_467 = 12'hf14 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_469 = 12'h300 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_471 = 12'h301 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_473 = 12'h302 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_475 = 12'h303 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_477 = 12'h304 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_479 = 12'h305 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_481 = 12'h306 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_483 = 12'h340 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_485 = 12'h341 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_487 = 12'h342 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_489 = 12'h343 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_491 = 12'h344 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_493 = 12'h3a0 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_495 = 12'h3a1 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_497 = 12'h3a2 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_499 = 12'h3a3 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_501 = 12'h3b0 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_503 = 12'h3b1 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_505 = 12'h3b2 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_507 = 12'h3b3 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_509 = 12'h3b4 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_511 = 12'h3b5 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_513 = 12'h3b6 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_515 = 12'h3b7 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_517 = 12'h3b8 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_519 = 12'h3b9 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_521 = 12'h3ba == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_523 = 12'h3bb == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_525 = 12'h3bc == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_527 = 12'h3bd == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_529 = 12'h3be == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_531 = 12'h3bf == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_533 = 12'hb00 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_535 = 12'hb02 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_537 = 12'hb80 == io_write_addr; // @[Lookup.scala 31:38]
  wire  _T_539 = 12'hb82 == io_write_addr; // @[Lookup.scala 31:38]
  wire [31:0] _T_543 = _T_539 ? minstret_data[63:32] : 32'h0; // @[Lookup.scala 33:37]
  wire [31:0] _T_544 = _T_537 ? mcycle_data[63:32] : _T_543; // @[Lookup.scala 33:37]
  wire [31:0] _T_545 = _T_535 ? minstret_data[31:0] : _T_544; // @[Lookup.scala 33:37]
  wire [31:0] _T_546 = _T_533 ? mcycle_data[31:0] : _T_545; // @[Lookup.scala 33:37]
  wire [31:0] _T_547 = _T_531 ? 32'h0 : _T_546; // @[Lookup.scala 33:37]
  wire [31:0] _T_548 = _T_529 ? 32'h0 : _T_547; // @[Lookup.scala 33:37]
  wire [31:0] _T_549 = _T_527 ? 32'h0 : _T_548; // @[Lookup.scala 33:37]
  wire [31:0] _T_550 = _T_525 ? 32'h0 : _T_549; // @[Lookup.scala 33:37]
  wire [31:0] _T_551 = _T_523 ? 32'h0 : _T_550; // @[Lookup.scala 33:37]
  wire [31:0] _T_552 = _T_521 ? 32'h0 : _T_551; // @[Lookup.scala 33:37]
  wire [31:0] _T_553 = _T_519 ? 32'h0 : _T_552; // @[Lookup.scala 33:37]
  wire [31:0] _T_554 = _T_517 ? 32'h0 : _T_553; // @[Lookup.scala 33:37]
  wire [31:0] _T_555 = _T_515 ? 32'h0 : _T_554; // @[Lookup.scala 33:37]
  wire [31:0] _T_556 = _T_513 ? 32'h0 : _T_555; // @[Lookup.scala 33:37]
  wire [31:0] _T_557 = _T_511 ? 32'h0 : _T_556; // @[Lookup.scala 33:37]
  wire [31:0] _T_558 = _T_509 ? 32'h0 : _T_557; // @[Lookup.scala 33:37]
  wire [31:0] _T_559 = _T_507 ? 32'h0 : _T_558; // @[Lookup.scala 33:37]
  wire [31:0] _T_560 = _T_505 ? 32'h0 : _T_559; // @[Lookup.scala 33:37]
  wire [31:0] _T_561 = _T_503 ? 32'h0 : _T_560; // @[Lookup.scala 33:37]
  wire [31:0] _T_562 = _T_501 ? 32'h0 : _T_561; // @[Lookup.scala 33:37]
  wire [31:0] _T_563 = _T_499 ? 32'h0 : _T_562; // @[Lookup.scala 33:37]
  wire [31:0] _T_564 = _T_497 ? 32'h0 : _T_563; // @[Lookup.scala 33:37]
  wire [31:0] _T_565 = _T_495 ? 32'h0 : _T_564; // @[Lookup.scala 33:37]
  wire [31:0] _T_566 = _T_493 ? 32'h0 : _T_565; // @[Lookup.scala 33:37]
  wire [31:0] _T_567 = _T_491 ? _T_142 : _T_566; // @[Lookup.scala 33:37]
  wire [31:0] _T_568 = _T_489 ? mtval_data : _T_567; // @[Lookup.scala 33:37]
  wire [31:0] _T_569 = _T_487 ? _T_130 : _T_568; // @[Lookup.scala 33:37]
  wire [31:0] _T_570 = _T_485 ? mepc_data : _T_569; // @[Lookup.scala 33:37]
  wire [31:0] _T_571 = _T_483 ? mscratch_data : _T_570; // @[Lookup.scala 33:37]
  wire [31:0] _T_572 = _T_481 ? 32'h0 : _T_571; // @[Lookup.scala 33:37]
  wire [31:0] _T_573 = _T_479 ? _T_129 : _T_572; // @[Lookup.scala 33:37]
  wire [31:0] _T_574 = _T_477 ? _T_47 : _T_573; // @[Lookup.scala 33:37]
  wire [31:0] _T_575 = _T_475 ? mideleg_data : _T_574; // @[Lookup.scala 33:37]
  wire [31:0] _T_576 = _T_473 ? medeleg_data : _T_575; // @[Lookup.scala 33:37]
  wire [31:0] _T_577 = _T_471 ? 32'h40141101 : _T_576; // @[Lookup.scala 33:37]
  wire [31:0] _T_578 = _T_469 ? _T_31 : _T_577; // @[Lookup.scala 33:37]
  wire [31:0] _T_579 = _T_467 ? 32'h0 : _T_578; // @[Lookup.scala 33:37]
  wire [31:0] _T_580 = _T_465 ? 32'h0 : _T_579; // @[Lookup.scala 33:37]
  wire [31:0] _T_581 = _T_463 ? 32'h0 : _T_580; // @[Lookup.scala 33:37]
  wire [31:0] _T_582 = _T_461 ? 32'h0 : _T_581; // @[Lookup.scala 33:37]
  wire [31:0] _T_583 = _T_459 ? _T_94 : _T_582; // @[Lookup.scala 33:37]
  wire [31:0] _T_584 = _T_457 ? _T_92 : _T_583; // @[Lookup.scala 33:37]
  wire [31:0] _T_585 = _T_455 ? stval_data : _T_584; // @[Lookup.scala 33:37]
  wire [31:0] _T_586 = _T_453 ? _T_84 : _T_585; // @[Lookup.scala 33:37]
  wire [31:0] _T_587 = _T_451 ? sepc_data : _T_586; // @[Lookup.scala 33:37]
  wire [31:0] _T_588 = _T_449 ? sscratch_data : _T_587; // @[Lookup.scala 33:37]
  wire [31:0] _T_589 = _T_447 ? 32'h0 : _T_588; // @[Lookup.scala 33:37]
  wire [31:0] _T_590 = _T_445 ? _T_83 : _T_589; // @[Lookup.scala 33:37]
  wire [31:0] _T_591 = _T_443 ? _T_82 : _T_590; // @[Lookup.scala 33:37]
  wire [31:0] _T_592 = _T_441 ? _T_74 : _T_591; // @[Lookup.scala 33:37]
  wire [31:0] _T_593 = _T_439 ? minstret_data[63:32] : _T_592; // @[Lookup.scala 33:37]
  wire [31:0] _T_594 = _T_437 ? mcycle_data[63:32] : _T_593; // @[Lookup.scala 33:37]
  wire [31:0] _T_595 = _T_435 ? minstret_data[31:0] : _T_594; // @[Lookup.scala 33:37]
  wire [31:0] csrData = _T_433 ? mcycle_data[31:0] : _T_595; // @[Lookup.scala 33:37]
  wire  _T_706 = io_write_op != 3'h0; // @[CsrFile.scala 148:31]
  wire  _T_707 = io_write_op != 3'h1; // @[CsrFile.scala 148:58]
  wire  writeEn = _T_706 & _T_707; // @[CsrFile.scala 148:43]
  wire [31:0] _T_708 = csrData | io_write_data; // @[CsrFile.scala 152:25]
  wire [31:0] _T_709 = ~io_write_data; // @[CsrFile.scala 153:27]
  wire [31:0] _T_710 = csrData & _T_709; // @[CsrFile.scala 153:25]
  wire  _T_711 = 3'h5 == io_write_op; // @[Mux.scala 68:19]
  wire [31:0] _T_712 = _T_711 ? _T_710 : 32'h0; // @[Mux.scala 68:16]
  wire  _T_713 = 3'h4 == io_write_op; // @[Mux.scala 68:19]
  wire [31:0] _T_714 = _T_713 ? _T_708 : _T_712; // @[Mux.scala 68:16]
  wire  _T_715 = 3'h3 == io_write_op; // @[Mux.scala 68:19]
  wire [31:0] _T_716 = _T_715 ? io_write_data : _T_714; // @[Mux.scala 68:16]
  wire  _T_717 = 3'h2 == io_write_op; // @[Mux.scala 68:19]
  wire [31:0] writeData = _T_717 ? io_write_data : _T_716; // @[Mux.scala 68:16]
  wire [31:0] flagIntS = _T_92 & _T_82; // @[CsrFile.scala 157:30]
  wire [31:0] flagIntM = _T_142 & _T_47; // @[CsrFile.scala 158:30]
  wire  _T_758 = mode < 2'h1; // @[CsrFile.scala 159:28]
  wire  _T_759 = mode == 2'h1; // @[CsrFile.scala 160:33]
  wire  _T_760 = _T_759 & mstatus_sie; // @[CsrFile.scala 160:48]
  wire  _T_761 = _T_758 | _T_760; // @[CsrFile.scala 159:41]
  wire [31:0] _T_762 = flagIntS & mideleg_data; // @[CsrFile.scala 161:33]
  wire  _T_763 = _T_762 != 32'h0; // @[CsrFile.scala 161:51]
  wire  hasIntS = _T_761 & _T_763; // @[CsrFile.scala 159:22]
  wire  _T_764 = mode <= 2'h1; // @[CsrFile.scala 162:28]
  wire  _T_765 = _T_764 | mstatus_mie; // @[CsrFile.scala 162:42]
  wire [31:0] _T_766 = ~mideleg_data; // @[CsrFile.scala 163:35]
  wire [31:0] _T_767 = flagIntM & _T_766; // @[CsrFile.scala 163:33]
  wire  _T_768 = _T_767 != 32'h0; // @[CsrFile.scala 163:52]
  wire  hasIntM = _T_765 & _T_768; // @[CsrFile.scala 162:22]
  wire  hasInt = hasIntM | hasIntS; // @[CsrFile.scala 164:27]
  wire  _T_769 = ~hasIntM; // @[CsrFile.scala 165:29]
  wire  handIntS = hasInt & _T_769; // @[CsrFile.scala 165:26]
  wire  _T_770 = ~hasInt; // @[CsrFile.scala 166:40]
  wire  hasExc = io_except_hasTrap & _T_770; // @[CsrFile.scala 166:37]
  wire [31:0] _T_772 = medeleg_data >> io_except_excCause[4:0]; // @[CsrFile.scala 167:45]
  wire  hasExcS = hasExc & _T_772[0]; // @[CsrFile.scala 167:26]
  wire  _T_775 = ~mode[1]; // @[CsrFile.scala 168:19]
  wire  handExcS = _T_775 & hasExcS; // @[CsrFile.scala 168:28]
  wire [31:0] _T_776 = {{9'd0}, flagIntS[31:9]}; // @[CsrFile.scala 169:31]
  wire [31:0] _T_778 = {{1'd0}, flagIntS[31:1]}; // @[CsrFile.scala 170:31]
  wire [30:0] _T_780 = _T_778[0] ? 31'h1 : 31'h5; // @[CsrFile.scala 170:22]
  wire [30:0] intCauseS = _T_776[0] ? 31'h9 : _T_780; // @[CsrFile.scala 169:22]
  wire [31:0] _T_781 = {{11'd0}, flagIntM[31:11]}; // @[CsrFile.scala 172:31]
  wire [31:0] _T_783 = {{3'd0}, flagIntM[31:3]}; // @[CsrFile.scala 173:31]
  wire [31:0] _T_785 = {{7'd0}, flagIntM[31:7]}; // @[CsrFile.scala 174:31]
  wire [30:0] _T_787 = _T_785[0] ? 31'h7 : intCauseS; // @[CsrFile.scala 174:22]
  wire [30:0] _T_788 = _T_783[0] ? 31'h3 : _T_787; // @[CsrFile.scala 173:22]
  wire [30:0] intCauseM = _T_781[0] ? 31'hb : _T_788; // @[CsrFile.scala 172:22]
  wire [30:0] intCause = handIntS ? intCauseS : intCauseM; // @[CsrFile.scala 176:22]
  wire [31:0] _T_789 = {1'h1,intCause}; // @[Cat.scala 30:58]
  wire [31:0] _T_790 = {1'h0,io_except_excCause}; // @[Cat.scala 30:58]
  wire [31:0] cause = hasInt ? _T_789 : _T_790; // @[CsrFile.scala 177:22]
  wire  _T_792 = stvec_mode[0] & hasInt; // @[CsrFile.scala 179:37]
  wire [29:0] _T_795 = stvec_base + cause[29:0]; // @[CsrFile.scala 179:60]
  wire [29:0] _T_796 = _T_792 ? _T_795 : stvec_base; // @[CsrFile.scala 179:22]
  wire [31:0] trapVecS = {_T_796, 2'h0}; // @[CsrFile.scala 180:35]
  wire  _T_798 = mtvec_mode[0] & hasInt; // @[CsrFile.scala 181:37]
  wire [29:0] _T_801 = mtvec_base + cause[29:0]; // @[CsrFile.scala 181:60]
  wire [29:0] _T_802 = _T_798 ? _T_801 : mtvec_base; // @[CsrFile.scala 181:22]
  wire [31:0] trapVecM = {_T_802, 2'h0}; // @[CsrFile.scala 182:35]
  wire  _T_803 = handIntS | handExcS; // @[CsrFile.scala 183:32]
  wire [1:0] sretMode = {1'h0,sstatus_spp}; // @[Cat.scala 30:58]
  wire  _T_812 = ~writeEn; // @[CsrFile.scala 204:44]
  wire  _T_813 = io_except_hasTrap & _T_812; // @[CsrFile.scala 204:41]
  wire [63:0] _T_815 = mcycle_data + 64'h1; // @[CsrFile.scala 208:30]
  wire [63:0] _T_817 = minstret_data + 64'h1; // @[CsrFile.scala 210:36]
  wire  _T_818 = io_write_addr == 12'h100; // @[CsrFile.scala 218:25]
  wire [8:0] _T_865 = {writeData[8],_T_31[7:6],writeData[5],_T_31[4],_T_31[3:2],writeData[1],_T_31[0]}; // @[CSR.scala 21:18]
  wire [31:0] _T_873 = {_T_31[31],_T_31[30:20],_T_31[19],writeData[18],_T_31[17],_T_31[16:15],_T_31[14:13],_T_31[12:9],_T_865}; // @[CSR.scala 21:18]
  wire  _T_881 = io_write_addr == 12'h104; // @[CsrFile.scala 221:25]
  wire [31:0] _T_915 = {_T_47[31:10],writeData[9],_T_47[8],_T_47[7:6],writeData[5],_T_47[4],_T_47[3:2],writeData[1],_T_47[0]}; // @[CSR.scala 21:18]
  wire  _T_922 = io_write_addr == 12'h144; // @[CsrFile.scala 224:25]
  wire [31:0] _T_935 = {21'h0,1'h0,mipReal_seip,3'h0,mipReal_stip,1'h0,1'h0,1'h0,mipReal_ssip,1'h0}; // @[CSR.scala 19:24]
  wire [31:0] _T_954 = {_T_935[31:10],_T_935[9],_T_935[8],_T_935[7:6],_T_935[5],_T_935[4],_T_935[3:2],writeData[1],_T_935[0]}; // @[CSR.scala 21:18]
  wire  _T_958 = io_write_addr == 12'hb00; // @[CsrFile.scala 227:25]
  wire [63:0] _T_960 = {mcycle_data[63:32],writeData}; // @[Cat.scala 30:58]
  wire  _T_961 = io_write_addr == 12'hb02; // @[CsrFile.scala 230:25]
  wire [63:0] _T_963 = {minstret_data[63:32],writeData}; // @[Cat.scala 30:58]
  wire  _T_964 = io_write_addr == 12'hb80; // @[CsrFile.scala 233:25]
  wire [63:0] _T_966 = {writeData,mcycle_data[31:0]}; // @[Cat.scala 30:58]
  wire  _T_967 = io_write_addr == 12'hb82; // @[CsrFile.scala 236:25]
  wire [63:0] _T_969 = {writeData,minstret_data[31:0]}; // @[Cat.scala 30:58]
  wire  _T_970 = io_write_addr == 12'h105; // @[CsrFile.scala 239:25]
  wire  _T_973 = io_write_addr == 12'h140; // @[CsrFile.scala 240:25]
  wire  _T_977 = io_write_addr == 12'h141; // @[CsrFile.scala 241:25]
  wire [31:0] _T_979 = {writeData[31:2],2'h0}; // @[Cat.scala 30:58]
  wire  _T_980 = io_write_addr == 12'h142; // @[CsrFile.scala 242:25]
  wire  _T_983 = io_write_addr == 12'h143; // @[CsrFile.scala 243:25]
  wire  _T_987 = io_write_addr == 12'h180; // @[CsrFile.scala 244:25]
  wire  _T_990 = io_write_addr == 12'h300; // @[CsrFile.scala 245:25]
  wire  _T_998 = io_write_addr == 12'h302; // @[CsrFile.scala 246:25]
  wire [6:0] _T_1008 = {writeData[6],1'h0,writeData[4:2],1'h0,writeData[0]}; // @[Cat.scala 30:58]
  wire [15:0] _T_1014 = {writeData[15],1'h0,writeData[13:12],2'h0,writeData[9:8],1'h0,_T_1008}; // @[Cat.scala 30:58]
  wire  _T_1015 = io_write_addr == 12'h303; // @[CsrFile.scala 247:25]
  wire [11:0] _T_1024 = {2'h0,writeData[9],3'h0,writeData[5],3'h0,writeData[1],1'h0}; // @[Cat.scala 30:58]
  wire  _T_1025 = io_write_addr == 12'h304; // @[CsrFile.scala 248:25]
  wire  _T_1032 = io_write_addr == 12'h305; // @[CsrFile.scala 249:25]
  wire  _T_1035 = io_write_addr == 12'h340; // @[CsrFile.scala 250:25]
  wire  _T_1039 = io_write_addr == 12'h341; // @[CsrFile.scala 251:25]
  wire  _T_1042 = io_write_addr == 12'h342; // @[CsrFile.scala 252:25]
  wire  _T_1045 = io_write_addr == 12'h343; // @[CsrFile.scala 253:25]
  wire  _T_1049 = io_write_addr == 12'h344; // @[CsrFile.scala 254:25]
  wire [31:0] _T_1055 = {io_except_excPc[31:2],2'h0}; // @[Cat.scala 30:58]
  wire  _GEN_59 = _T_803 ? mstatus_sie : mstatus_spie; // @[CsrFile.scala 268:40]
  wire  _GEN_66 = _T_803 ? mstatus_mpie : mstatus_mie; // @[CsrFile.scala 268:40]
  wire  _GEN_67 = _T_803 & mstatus_mie; // @[CsrFile.scala 268:40]
  wire  _GEN_70 = io_except_isMret | _GEN_66; // @[CsrFile.scala 263:36]
  wire  _GEN_76 = io_except_isMret ? mstatus_spie : _GEN_59; // @[CsrFile.scala 263:36]
  wire  _GEN_84 = io_except_isSret | _GEN_76; // @[CsrFile.scala 257:29]
  assign io_read_valid = readValid & modeValid; // @[CsrFile.scala 289:17]
  assign io_read_data = _T_148 ? mcycle_data[31:0] : _T_310; // @[CsrFile.scala 290:17]
  assign io_hasInt = hasIntM | hasIntS; // @[CsrFile.scala 293:15]
  assign io_busy = _T_706 & _T_707; // @[CsrFile.scala 294:15]
  assign io_mode = mode; // @[CsrFile.scala 295:15]
  assign io_sepc = sepc_data; // @[CsrFile.scala 296:15]
  assign io_mepc = mepc_data; // @[CsrFile.scala 297:15]
  assign io_trapVec = _T_803 ? trapVecS : trapVecM; // @[CsrFile.scala 298:15]
  assign io_pageEn = _T_775 & satp_mode; // @[CsrFile.scala 301:15]
  assign io_basePpn = satp_ppn; // @[CsrFile.scala 302:15]
  assign io_sum = mstatus_sum; // @[CsrFile.scala 303:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mode = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mstatus_sum = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mstatus_mpp = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  mstatus_spp = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mstatus_mpie = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mstatus_spie = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  mstatus_mie = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mstatus_sie = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  medeleg_data = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  mideleg_data = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mie_meie = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mie_seie = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  mie_mtie = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  mie_stie = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  mie_msie = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  mie_ssie = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  mtvec_base = _RAND_16[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  mtvec_mode = _RAND_17[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  mscratch_data = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  mepc_data = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  mcause_int = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  mcause_code = _RAND_21[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mtval_data = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mipReal_seip = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  mipReal_stip = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mipReal_ssip = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {2{`RANDOM}};
  mcycle_data = _RAND_26[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  minstret_data = _RAND_27[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  stvec_base = _RAND_28[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  stvec_mode = _RAND_29[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  sscratch_data = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  sepc_data = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  scause_int = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  scause_code = _RAND_33[30:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  stval_data = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  satp_mode = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  satp_ppn = _RAND_36[21:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      mode <= 2'h3;
    end else if (_T_813) begin
      if (hasInt) begin
        if (handIntS) begin
          mode <= 2'h1;
        end else begin
          mode <= 2'h3;
        end
      end else if (io_except_isSret) begin
        mode <= sretMode;
      end else if (io_except_isMret) begin
        mode <= mstatus_mpp;
      end else if (handExcS) begin
        mode <= 2'h1;
      end else begin
        mode <= 2'h3;
      end
    end
    if (reset) begin
      mstatus_sum <= 1'h0;
    end else if (writeEn) begin
      if (_T_990) begin
        mstatus_sum <= writeData[18];
      end else if (_T_818) begin
        mstatus_sum <= _T_873[18];
      end
    end
    if (reset) begin
      mstatus_mpp <= 2'h0;
    end else if (writeEn) begin
      if (_T_990) begin
        mstatus_mpp <= writeData[12:11];
      end else if (_T_818) begin
        mstatus_mpp <= _T_873[12:11];
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        if (io_except_isMret) begin
          mstatus_mpp <= 2'h0;
        end else if (!(_T_803)) begin
          mstatus_mpp <= mode;
        end
      end
    end
    if (reset) begin
      mstatus_spp <= 1'h0;
    end else if (writeEn) begin
      if (_T_990) begin
        mstatus_spp <= writeData[8];
      end else if (_T_818) begin
        mstatus_spp <= _T_873[8];
      end
    end else if (io_except_hasTrap) begin
      if (io_except_isSret) begin
        mstatus_spp <= 1'h0;
      end else if (!(io_except_isMret)) begin
        if (_T_803) begin
          mstatus_spp <= mode[0];
        end
      end
    end
    if (reset) begin
      mstatus_mpie <= 1'h0;
    end else if (writeEn) begin
      if (_T_990) begin
        mstatus_mpie <= writeData[7];
      end else if (_T_818) begin
        mstatus_mpie <= _T_873[7];
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        mstatus_mpie <= _GEN_70;
      end
    end
    if (reset) begin
      mstatus_spie <= 1'h0;
    end else if (writeEn) begin
      if (_T_990) begin
        mstatus_spie <= writeData[5];
      end else if (_T_818) begin
        mstatus_spie <= _T_873[5];
      end
    end else if (io_except_hasTrap) begin
      mstatus_spie <= _GEN_84;
    end
    if (reset) begin
      mstatus_mie <= 1'h0;
    end else if (writeEn) begin
      if (_T_990) begin
        mstatus_mie <= writeData[3];
      end else if (_T_818) begin
        mstatus_mie <= _T_873[3];
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        if (io_except_isMret) begin
          mstatus_mie <= mstatus_mpie;
        end else begin
          mstatus_mie <= _GEN_67;
        end
      end
    end
    if (reset) begin
      mstatus_sie <= 1'h0;
    end else if (writeEn) begin
      if (_T_990) begin
        mstatus_sie <= writeData[1];
      end else if (_T_818) begin
        mstatus_sie <= _T_873[1];
      end
    end else if (io_except_hasTrap) begin
      if (io_except_isSret) begin
        mstatus_sie <= mstatus_spie;
      end else if (!(io_except_isMret)) begin
        if (_T_803) begin
          mstatus_sie <= 1'h0;
        end
      end
    end
    if (reset) begin
      medeleg_data <= 32'h0;
    end else if (writeEn) begin
      if (_T_998) begin
        medeleg_data <= {{16'd0}, _T_1014};
      end
    end
    if (reset) begin
      mideleg_data <= 32'h0;
    end else if (writeEn) begin
      if (_T_1015) begin
        mideleg_data <= {{20'd0}, _T_1024};
      end
    end
    if (reset) begin
      mie_meie <= 1'h0;
    end else if (writeEn) begin
      if (_T_1025) begin
        mie_meie <= writeData[11];
      end else if (_T_881) begin
        mie_meie <= _T_915[11];
      end
    end
    if (reset) begin
      mie_seie <= 1'h0;
    end else if (writeEn) begin
      if (_T_1025) begin
        mie_seie <= writeData[9];
      end else if (_T_881) begin
        mie_seie <= _T_915[9];
      end
    end
    if (reset) begin
      mie_mtie <= 1'h0;
    end else if (writeEn) begin
      if (_T_1025) begin
        mie_mtie <= writeData[7];
      end else if (_T_881) begin
        mie_mtie <= _T_915[7];
      end
    end
    if (reset) begin
      mie_stie <= 1'h0;
    end else if (writeEn) begin
      if (_T_1025) begin
        mie_stie <= writeData[5];
      end else if (_T_881) begin
        mie_stie <= _T_915[5];
      end
    end
    if (reset) begin
      mie_msie <= 1'h0;
    end else if (writeEn) begin
      if (_T_1025) begin
        mie_msie <= writeData[3];
      end else if (_T_881) begin
        mie_msie <= _T_915[3];
      end
    end
    if (reset) begin
      mie_ssie <= 1'h0;
    end else if (writeEn) begin
      if (_T_1025) begin
        mie_ssie <= writeData[1];
      end else if (_T_881) begin
        mie_ssie <= _T_915[1];
      end
    end
    if (reset) begin
      mtvec_base <= 30'h0;
    end else if (writeEn) begin
      if (_T_1032) begin
        mtvec_base <= writeData[31:2];
      end
    end
    if (reset) begin
      mtvec_mode <= 2'h0;
    end else if (writeEn) begin
      if (_T_1032) begin
        mtvec_mode <= {{1'd0}, writeData[0]};
      end
    end
    if (reset) begin
      mscratch_data <= 32'h0;
    end else if (writeEn) begin
      if (_T_1035) begin
        if (_T_717) begin
          mscratch_data <= io_write_data;
        end else if (_T_715) begin
          mscratch_data <= io_write_data;
        end else if (_T_713) begin
          mscratch_data <= _T_708;
        end else if (_T_711) begin
          mscratch_data <= _T_710;
        end else begin
          mscratch_data <= 32'h0;
        end
      end
    end
    if (reset) begin
      mepc_data <= 32'h0;
    end else if (writeEn) begin
      if (_T_1039) begin
        mepc_data <= _T_979;
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        if (!(io_except_isMret)) begin
          if (!(_T_803)) begin
            mepc_data <= _T_1055;
          end
        end
      end
    end
    if (reset) begin
      mcause_int <= 1'h0;
    end else if (writeEn) begin
      if (_T_1042) begin
        mcause_int <= writeData[31];
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        if (!(io_except_isMret)) begin
          if (!(_T_803)) begin
            mcause_int <= cause[31];
          end
        end
      end
    end
    if (reset) begin
      mcause_code <= 31'h0;
    end else if (writeEn) begin
      if (_T_1042) begin
        mcause_code <= {{27'd0}, writeData[3:0]};
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        if (!(io_except_isMret)) begin
          if (!(_T_803)) begin
            mcause_code <= {{27'd0}, cause[3:0]};
          end
        end
      end
    end
    if (reset) begin
      mtval_data <= 32'h0;
    end else if (writeEn) begin
      if (_T_1045) begin
        if (_T_717) begin
          mtval_data <= io_write_data;
        end else if (_T_715) begin
          mtval_data <= io_write_data;
        end else if (_T_713) begin
          mtval_data <= _T_708;
        end else if (_T_711) begin
          mtval_data <= _T_710;
        end else begin
          mtval_data <= 32'h0;
        end
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        if (!(io_except_isMret)) begin
          if (!(_T_803)) begin
            mtval_data <= io_except_excValue;
          end
        end
      end
    end
    if (reset) begin
      mipReal_seip <= 1'h0;
    end else if (writeEn) begin
      if (_T_1049) begin
        mipReal_seip <= writeData[9];
      end else if (_T_922) begin
        mipReal_seip <= _T_954[9];
      end
    end
    if (reset) begin
      mipReal_stip <= 1'h0;
    end else if (writeEn) begin
      if (_T_1049) begin
        mipReal_stip <= writeData[5];
      end else if (_T_922) begin
        mipReal_stip <= _T_954[5];
      end
    end
    if (reset) begin
      mipReal_ssip <= 1'h0;
    end else if (writeEn) begin
      if (_T_1049) begin
        mipReal_ssip <= writeData[1];
      end else if (_T_922) begin
        mipReal_ssip <= _T_954[1];
      end
    end
    if (reset) begin
      mcycle_data <= 64'h0;
    end else if (writeEn) begin
      if (_T_964) begin
        mcycle_data <= _T_966;
      end else if (_T_958) begin
        mcycle_data <= _T_960;
      end else begin
        mcycle_data <= _T_815;
      end
    end else begin
      mcycle_data <= _T_815;
    end
    if (reset) begin
      minstret_data <= 64'h0;
    end else if (writeEn) begin
      if (_T_967) begin
        minstret_data <= _T_969;
      end else if (_T_961) begin
        minstret_data <= _T_963;
      end else if (io_write_retired) begin
        minstret_data <= _T_817;
      end
    end else if (io_write_retired) begin
      minstret_data <= _T_817;
    end
    if (reset) begin
      stvec_base <= 30'h0;
    end else if (writeEn) begin
      if (_T_970) begin
        stvec_base <= writeData[31:2];
      end
    end
    if (reset) begin
      stvec_mode <= 2'h0;
    end else if (writeEn) begin
      if (_T_970) begin
        stvec_mode <= {{1'd0}, writeData[0]};
      end
    end
    if (reset) begin
      sscratch_data <= 32'h0;
    end else if (writeEn) begin
      if (_T_973) begin
        if (_T_717) begin
          sscratch_data <= io_write_data;
        end else if (_T_715) begin
          sscratch_data <= io_write_data;
        end else if (_T_713) begin
          sscratch_data <= _T_708;
        end else if (_T_711) begin
          sscratch_data <= _T_710;
        end else begin
          sscratch_data <= 32'h0;
        end
      end
    end
    if (reset) begin
      sepc_data <= 32'h0;
    end else if (writeEn) begin
      if (_T_977) begin
        sepc_data <= _T_979;
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        if (!(io_except_isMret)) begin
          if (_T_803) begin
            sepc_data <= _T_1055;
          end
        end
      end
    end
    if (reset) begin
      scause_int <= 1'h0;
    end else if (writeEn) begin
      if (_T_980) begin
        scause_int <= writeData[31];
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        if (!(io_except_isMret)) begin
          if (_T_803) begin
            scause_int <= cause[31];
          end
        end
      end
    end
    if (reset) begin
      scause_code <= 31'h0;
    end else if (writeEn) begin
      if (_T_980) begin
        scause_code <= {{27'd0}, writeData[3:0]};
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        if (!(io_except_isMret)) begin
          if (_T_803) begin
            scause_code <= {{27'd0}, cause[3:0]};
          end
        end
      end
    end
    if (reset) begin
      stval_data <= 32'h0;
    end else if (writeEn) begin
      if (_T_983) begin
        if (_T_717) begin
          stval_data <= io_write_data;
        end else if (_T_715) begin
          stval_data <= io_write_data;
        end else if (_T_713) begin
          stval_data <= _T_708;
        end else if (_T_711) begin
          stval_data <= _T_710;
        end else begin
          stval_data <= 32'h0;
        end
      end
    end else if (io_except_hasTrap) begin
      if (!(io_except_isSret)) begin
        if (!(io_except_isMret)) begin
          if (_T_803) begin
            stval_data <= io_except_excValue;
          end
        end
      end
    end
    if (reset) begin
      satp_mode <= 1'h0;
    end else if (writeEn) begin
      if (_T_987) begin
        satp_mode <= writeData[31];
      end
    end
    if (reset) begin
      satp_ppn <= 22'h0;
    end else if (writeEn) begin
      if (_T_987) begin
        satp_ppn <= writeData[21:0];
      end
    end
  end
endmodule
module ExclusiveMonitor(
  input         clock,
  input         reset,
  input         io_flush,
  input  [31:0] io_check_addr,
  output        io_check_valid,
  input  [31:0] io_update_addr,
  input         io_update_set,
  input         io_update_clear
);
  reg  flag; // @[ExclusiveMonitor.scala 20:22]
  reg [31:0] _RAND_0;
  reg [31:0] addr; // @[ExclusiveMonitor.scala 21:22]
  reg [31:0] _RAND_1;
  wire  _T = io_update_addr == addr; // @[ExclusiveMonitor.scala 23:56]
  wire  _T_1 = io_update_clear & _T; // @[ExclusiveMonitor.scala 23:38]
  wire  _T_2 = io_flush | _T_1; // @[ExclusiveMonitor.scala 23:18]
  wire  _GEN_0 = io_update_set | flag; // @[ExclusiveMonitor.scala 26:31]
  wire  _T_3 = addr == io_check_addr; // @[ExclusiveMonitor.scala 31:34]
  assign io_check_valid = flag & _T_3; // @[ExclusiveMonitor.scala 31:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  flag = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  addr = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      flag <= 1'h0;
    end else if (_T_2) begin
      flag <= 1'h0;
    end else begin
      flag <= _GEN_0;
    end
    if (reset) begin
      addr <= 32'h0;
    end else if (_T_2) begin
      addr <= 32'h0;
    end else if (io_update_set) begin
      addr <= io_update_addr;
    end
  end
endmodule
module HazardResolver(
  input         io_regRead1_en,
  input  [4:0]  io_regRead1_addr,
  output [31:0] io_regRead1_data,
  input         io_regRead2_en,
  input  [4:0]  io_regRead2_addr,
  output [31:0] io_regRead2_data,
  input  [2:0]  io_csrRead_op,
  output        io_csrRead_valid,
  input  [11:0] io_csrRead_addr,
  output [31:0] io_csrRead_data,
  input  [31:0] io_check_addr,
  output        io_check_valid,
  input         io_aluReg_en,
  input  [4:0]  io_aluReg_addr,
  input  [31:0] io_aluReg_data,
  input         io_aluReg_load,
  input         io_memReg_en,
  input  [4:0]  io_memReg_addr,
  input  [31:0] io_memReg_data,
  input         io_memReg_load,
  input  [2:0]  io_memCsr_op,
  input  [11:0] io_memCsr_addr,
  input         io_wbReg_en,
  input  [4:0]  io_wbReg_addr,
  input  [31:0] io_wbReg_data,
  input  [2:0]  io_wbCsr_op,
  input  [11:0] io_wbCsr_addr,
  input  [31:0] io_wbExcMon_addr,
  input         io_wbExcMon_set,
  input         io_wbExcMon_clear,
  output        io_rf1_en,
  output [4:0]  io_rf1_addr,
  input  [31:0] io_rf1_data,
  output        io_rf2_en,
  output [4:0]  io_rf2_addr,
  input  [31:0] io_rf2_data,
  output [2:0]  io_csr_op,
  input         io_csr_valid,
  output [11:0] io_csr_addr,
  input  [31:0] io_csr_data,
  output [31:0] io_excMon_addr,
  input         io_excMon_valid,
  output        io_loadFlag,
  output        io_csrFlag
);
  wire  _T = io_regRead1_addr != 5'h0; // @[HazardResolver.scala 39:32]
  wire  _T_1 = io_regRead1_en & _T; // @[HazardResolver.scala 39:19]
  wire  _T_2 = io_regRead1_addr == io_aluReg_addr; // @[HazardResolver.scala 40:39]
  wire  _T_3 = io_aluReg_en & _T_2; // @[HazardResolver.scala 40:26]
  wire  _T_4 = io_regRead1_addr == io_memReg_addr; // @[HazardResolver.scala 42:46]
  wire  _T_5 = io_memReg_en & _T_4; // @[HazardResolver.scala 42:33]
  wire  _T_6 = io_regRead1_addr == io_wbReg_addr; // @[HazardResolver.scala 44:45]
  wire  _T_7 = io_wbReg_en & _T_6; // @[HazardResolver.scala 44:32]
  wire [31:0] _GEN_0 = _T_7 ? io_wbReg_data : io_rf1_data; // @[HazardResolver.scala 44:64]
  wire [31:0] _GEN_1 = _T_5 ? io_memReg_data : _GEN_0; // @[HazardResolver.scala 42:66]
  wire [31:0] _GEN_2 = _T_3 ? io_aluReg_data : _GEN_1; // @[HazardResolver.scala 40:59]
  wire  _T_8 = io_regRead2_addr != 5'h0; // @[HazardResolver.scala 39:32]
  wire  _T_9 = io_regRead2_en & _T_8; // @[HazardResolver.scala 39:19]
  wire  _T_10 = io_regRead2_addr == io_aluReg_addr; // @[HazardResolver.scala 40:39]
  wire  _T_11 = io_aluReg_en & _T_10; // @[HazardResolver.scala 40:26]
  wire  _T_12 = io_regRead2_addr == io_memReg_addr; // @[HazardResolver.scala 42:46]
  wire  _T_13 = io_memReg_en & _T_12; // @[HazardResolver.scala 42:33]
  wire  _T_14 = io_regRead2_addr == io_wbReg_addr; // @[HazardResolver.scala 44:45]
  wire  _T_15 = io_wbReg_en & _T_14; // @[HazardResolver.scala 44:32]
  wire [31:0] _GEN_4 = _T_15 ? io_wbReg_data : io_rf2_data; // @[HazardResolver.scala 44:64]
  wire [31:0] _GEN_5 = _T_13 ? io_memReg_data : _GEN_4; // @[HazardResolver.scala 42:66]
  wire [31:0] _GEN_6 = _T_11 ? io_aluReg_data : _GEN_5; // @[HazardResolver.scala 40:59]
  wire  _T_16 = io_wbExcMon_clear | io_wbExcMon_set; // @[HazardResolver.scala 55:29]
  wire  _T_17 = io_check_addr == io_wbExcMon_addr; // @[HazardResolver.scala 56:24]
  wire  _GEN_8 = io_wbExcMon_clear ? 1'h0 : 1'h1; // @[HazardResolver.scala 57:34]
  wire  _GEN_9 = _T_17 & _GEN_8; // @[HazardResolver.scala 56:46]
  wire  _T_19 = io_aluReg_load & _T_2; // @[HazardResolver.scala 71:34]
  wire  _T_21 = io_memReg_load & _T_4; // @[HazardResolver.scala 72:34]
  wire  _T_22 = _T_19 | _T_21; // @[HazardResolver.scala 73:25]
  wire  loadHazard1 = io_regRead1_en & _T_22; // @[HazardResolver.scala 73:13]
  wire  _T_24 = io_aluReg_load & _T_10; // @[HazardResolver.scala 71:34]
  wire  _T_26 = io_memReg_load & _T_12; // @[HazardResolver.scala 72:34]
  wire  _T_27 = _T_24 | _T_26; // @[HazardResolver.scala 73:25]
  wire  loadHazard2 = io_regRead2_en & _T_27; // @[HazardResolver.scala 73:13]
  wire  _T_28 = io_csrRead_op != 3'h0; // @[HazardResolver.scala 77:27]
  wire  _T_29 = io_csrRead_op != 3'h2; // @[HazardResolver.scala 77:50]
  wire  _T_30 = _T_28 & _T_29; // @[HazardResolver.scala 77:39]
  wire  _T_31 = io_memCsr_op != 3'h0; // @[HazardResolver.scala 78:32]
  wire  _T_32 = io_memCsr_op != 3'h1; // @[HazardResolver.scala 78:60]
  wire  _T_33 = _T_31 & _T_32; // @[HazardResolver.scala 78:44]
  wire  _T_34 = io_csrRead_addr == io_memCsr_addr; // @[HazardResolver.scala 79:29]
  wire  _T_35 = _T_33 & _T_34; // @[HazardResolver.scala 78:70]
  wire  _T_36 = io_wbCsr_op != 3'h0; // @[HazardResolver.scala 80:31]
  wire  _T_37 = io_wbCsr_op != 3'h1; // @[HazardResolver.scala 80:58]
  wire  _T_38 = _T_36 & _T_37; // @[HazardResolver.scala 80:43]
  wire  _T_39 = io_csrRead_addr == io_wbCsr_addr; // @[HazardResolver.scala 81:29]
  wire  _T_40 = _T_38 & _T_39; // @[HazardResolver.scala 80:68]
  wire  _T_41 = _T_35 | _T_40; // @[HazardResolver.scala 82:23]
  assign io_regRead1_data = _T_1 ? _GEN_2 : 32'h0; // @[HazardResolver.scala 41:19 HazardResolver.scala 43:19 HazardResolver.scala 45:19 HazardResolver.scala 47:19 HazardResolver.scala 50:17]
  assign io_regRead2_data = _T_9 ? _GEN_6 : 32'h0; // @[HazardResolver.scala 41:19 HazardResolver.scala 43:19 HazardResolver.scala 45:19 HazardResolver.scala 47:19 HazardResolver.scala 50:17]
  assign io_csrRead_valid = io_csr_valid; // @[HazardResolver.scala 104:10]
  assign io_csrRead_data = io_csr_data; // @[HazardResolver.scala 104:10]
  assign io_check_valid = _T_16 ? _GEN_9 : io_excMon_valid; // @[HazardResolver.scala 58:23 HazardResolver.scala 60:23 HazardResolver.scala 63:21 HazardResolver.scala 66:19]
  assign io_rf1_en = io_regRead1_en; // @[HazardResolver.scala 98:15]
  assign io_rf1_addr = io_regRead1_addr; // @[HazardResolver.scala 99:15]
  assign io_rf2_en = io_regRead2_en; // @[HazardResolver.scala 100:15]
  assign io_rf2_addr = io_regRead2_addr; // @[HazardResolver.scala 101:15]
  assign io_csr_op = io_csrRead_op; // @[HazardResolver.scala 104:10]
  assign io_csr_addr = io_csrRead_addr; // @[HazardResolver.scala 104:10]
  assign io_excMon_addr = io_check_addr; // @[HazardResolver.scala 107:19]
  assign io_loadFlag = loadHazard1 | loadHazard2; // @[HazardResolver.scala 110:15]
  assign io_csrFlag = _T_30 & _T_41; // @[HazardResolver.scala 111:15]
endmodule
module PipelineController(
  input         io_fetch,
  input         io_alu,
  input         io_mem,
  input         io_decFlush,
  input  [31:0] io_decTarget,
  input         io_memFlush,
  input  [31:0] io_memTarget,
  input         io_load,
  input         io_csr,
  input         io_except_hasTrap,
  input         io_except_isSret,
  input         io_except_isMret,
  input  [31:0] io_csrSepc,
  input  [31:0] io_csrMepc,
  input  [31:0] io_csrTvec,
  output        io_stallIf,
  output        io_stallId,
  output        io_stallEx,
  output        io_stallMm,
  output        io_stallWb,
  output        io_flush,
  output        io_flushIf,
  output [31:0] io_flushPc
);
  wire  _T = io_csr | io_alu; // @[PipelineController.scala 43:26]
  wire [4:0] _T_1 = io_fetch ? 5'h10 : 5'h0; // @[PipelineController.scala 45:18]
  wire [4:0] _T_2 = io_load ? 5'h18 : _T_1; // @[PipelineController.scala 44:18]
  wire [4:0] _T_3 = _T ? 5'h1c : _T_2; // @[PipelineController.scala 43:18]
  wire [4:0] stall = io_mem ? 5'h1e : _T_3; // @[PipelineController.scala 42:18]
  wire [31:0] _T_4 = io_except_isMret ? io_csrMepc : io_csrTvec; // @[PipelineController.scala 49:20]
  wire [31:0] excPc = io_except_isSret ? io_csrSepc : _T_4; // @[PipelineController.scala 48:20]
  wire  flushAll = io_except_hasTrap | io_memFlush; // @[PipelineController.scala 55:28]
  wire [31:0] _T_5 = io_memFlush ? io_memTarget : io_decTarget; // @[PipelineController.scala 58:22]
  assign io_stallIf = stall[4]; // @[PipelineController.scala 61:15]
  assign io_stallId = stall[3]; // @[PipelineController.scala 62:15]
  assign io_stallEx = stall[2]; // @[PipelineController.scala 63:15]
  assign io_stallMm = stall[1]; // @[PipelineController.scala 64:15]
  assign io_stallWb = stall[0]; // @[PipelineController.scala 65:15]
  assign io_flush = io_except_hasTrap | io_memFlush; // @[PipelineController.scala 68:15]
  assign io_flushIf = flushAll | io_decFlush; // @[PipelineController.scala 69:15]
  assign io_flushPc = io_except_hasTrap ? excPc : _T_5; // @[PipelineController.scala 70:15]
endmodule
module Core(
  input         clock,
  input         reset,
  input         io_irq_timer,
  input         io_irq_soft,
  input         io_irq_extern,
  output        io_tlb_en,
  output        io_tlb_flushInst,
  output        io_tlb_flushData,
  output [21:0] io_tlb_basePpn,
  output        io_tlb_sum,
  output        io_tlb_smode,
  output        io_cache_flushInst,
  output        io_cache_flushData,
  input         io_rom_valid,
  input         io_rom_fault,
  output [31:0] io_rom_addr,
  input  [31:0] io_rom_rdata,
  output        io_ram_en,
  input         io_ram_valid,
  input         io_ram_fault,
  output [3:0]  io_ram_wen,
  output [31:0] io_ram_addr,
  input  [31:0] io_ram_rdata,
  output [31:0] io_ram_wdata,
  output        io_debug_regWen,
  output [4:0]  io_debug_regWaddr,
  output [31:0] io_debug_regWdata,
  output [31:0] io_debug_pc
);
  wire  fetch_clock; // @[Core.scala 29:23]
  wire  fetch_reset; // @[Core.scala 29:23]
  wire  fetch_io_flush; // @[Core.scala 29:23]
  wire  fetch_io_stall; // @[Core.scala 29:23]
  wire  fetch_io_stallReq; // @[Core.scala 29:23]
  wire [31:0] fetch_io_flushPc; // @[Core.scala 29:23]
  wire  fetch_io_rom_valid; // @[Core.scala 29:23]
  wire  fetch_io_rom_fault; // @[Core.scala 29:23]
  wire [31:0] fetch_io_rom_addr; // @[Core.scala 29:23]
  wire  fetch_io_branch_branch; // @[Core.scala 29:23]
  wire  fetch_io_branch_jump; // @[Core.scala 29:23]
  wire  fetch_io_branch_taken; // @[Core.scala 29:23]
  wire [4:0] fetch_io_branch_index; // @[Core.scala 29:23]
  wire [31:0] fetch_io_branch_pc; // @[Core.scala 29:23]
  wire [31:0] fetch_io_branch_target; // @[Core.scala 29:23]
  wire  fetch_io_fetch_valid; // @[Core.scala 29:23]
  wire [31:0] fetch_io_fetch_pc; // @[Core.scala 29:23]
  wire  fetch_io_fetch_taken; // @[Core.scala 29:23]
  wire [31:0] fetch_io_fetch_target; // @[Core.scala 29:23]
  wire [4:0] fetch_io_fetch_predIndex; // @[Core.scala 29:23]
  wire  fetch_io_fetch_pageFault; // @[Core.scala 29:23]
  wire  ifid_clock; // @[Core.scala 30:23]
  wire  ifid_reset; // @[Core.scala 30:23]
  wire  ifid_io_flush; // @[Core.scala 30:23]
  wire  ifid_io_stallPrev; // @[Core.scala 30:23]
  wire  ifid_io_stallNext; // @[Core.scala 30:23]
  wire  ifid_io_prev_valid; // @[Core.scala 30:23]
  wire [31:0] ifid_io_prev_pc; // @[Core.scala 30:23]
  wire  ifid_io_prev_taken; // @[Core.scala 30:23]
  wire [31:0] ifid_io_prev_target; // @[Core.scala 30:23]
  wire [4:0] ifid_io_prev_predIndex; // @[Core.scala 30:23]
  wire  ifid_io_prev_pageFault; // @[Core.scala 30:23]
  wire  ifid_io_next_valid; // @[Core.scala 30:23]
  wire [31:0] ifid_io_next_pc; // @[Core.scala 30:23]
  wire  ifid_io_next_taken; // @[Core.scala 30:23]
  wire [31:0] ifid_io_next_target; // @[Core.scala 30:23]
  wire [4:0] ifid_io_next_predIndex; // @[Core.scala 30:23]
  wire  ifid_io_next_pageFault; // @[Core.scala 30:23]
  wire  decoder_clock; // @[Core.scala 31:23]
  wire  decoder_io_fetch_valid; // @[Core.scala 31:23]
  wire [31:0] decoder_io_fetch_pc; // @[Core.scala 31:23]
  wire  decoder_io_fetch_taken; // @[Core.scala 31:23]
  wire [31:0] decoder_io_fetch_target; // @[Core.scala 31:23]
  wire [4:0] decoder_io_fetch_predIndex; // @[Core.scala 31:23]
  wire  decoder_io_fetch_pageFault; // @[Core.scala 31:23]
  wire [31:0] decoder_io_inst; // @[Core.scala 31:23]
  wire  decoder_io_stallId; // @[Core.scala 31:23]
  wire  decoder_io_flushIf; // @[Core.scala 31:23]
  wire [31:0] decoder_io_flushPc; // @[Core.scala 31:23]
  wire  decoder_io_read1_en; // @[Core.scala 31:23]
  wire [4:0] decoder_io_read1_addr; // @[Core.scala 31:23]
  wire [31:0] decoder_io_read1_data; // @[Core.scala 31:23]
  wire  decoder_io_read2_en; // @[Core.scala 31:23]
  wire [4:0] decoder_io_read2_addr; // @[Core.scala 31:23]
  wire [31:0] decoder_io_read2_data; // @[Core.scala 31:23]
  wire  decoder_io_branch_branch; // @[Core.scala 31:23]
  wire  decoder_io_branch_jump; // @[Core.scala 31:23]
  wire  decoder_io_branch_taken; // @[Core.scala 31:23]
  wire [4:0] decoder_io_branch_index; // @[Core.scala 31:23]
  wire [31:0] decoder_io_branch_pc; // @[Core.scala 31:23]
  wire [31:0] decoder_io_branch_target; // @[Core.scala 31:23]
  wire [3:0] decoder_io_decoder_aluOp; // @[Core.scala 31:23]
  wire [31:0] decoder_io_decoder_opr1; // @[Core.scala 31:23]
  wire [31:0] decoder_io_decoder_opr2; // @[Core.scala 31:23]
  wire [3:0] decoder_io_decoder_mduOp; // @[Core.scala 31:23]
  wire [4:0] decoder_io_decoder_lsuOp; // @[Core.scala 31:23]
  wire [31:0] decoder_io_decoder_lsuData; // @[Core.scala 31:23]
  wire  decoder_io_decoder_regWen; // @[Core.scala 31:23]
  wire [4:0] decoder_io_decoder_regWaddr; // @[Core.scala 31:23]
  wire [2:0] decoder_io_decoder_csrOp; // @[Core.scala 31:23]
  wire [11:0] decoder_io_decoder_csrAddr; // @[Core.scala 31:23]
  wire [31:0] decoder_io_decoder_csrData; // @[Core.scala 31:23]
  wire [3:0] decoder_io_decoder_excType; // @[Core.scala 31:23]
  wire [31:0] decoder_io_decoder_excValue; // @[Core.scala 31:23]
  wire  decoder_io_decoder_valid; // @[Core.scala 31:23]
  wire [31:0] decoder_io_decoder_inst; // @[Core.scala 31:23]
  wire [31:0] decoder_io_decoder_currentPc; // @[Core.scala 31:23]
  wire  idex_clock; // @[Core.scala 32:23]
  wire  idex_reset; // @[Core.scala 32:23]
  wire  idex_io_flush; // @[Core.scala 32:23]
  wire  idex_io_stallPrev; // @[Core.scala 32:23]
  wire  idex_io_stallNext; // @[Core.scala 32:23]
  wire [3:0] idex_io_prev_aluOp; // @[Core.scala 32:23]
  wire [31:0] idex_io_prev_opr1; // @[Core.scala 32:23]
  wire [31:0] idex_io_prev_opr2; // @[Core.scala 32:23]
  wire [3:0] idex_io_prev_mduOp; // @[Core.scala 32:23]
  wire [4:0] idex_io_prev_lsuOp; // @[Core.scala 32:23]
  wire [31:0] idex_io_prev_lsuData; // @[Core.scala 32:23]
  wire  idex_io_prev_regWen; // @[Core.scala 32:23]
  wire [4:0] idex_io_prev_regWaddr; // @[Core.scala 32:23]
  wire [2:0] idex_io_prev_csrOp; // @[Core.scala 32:23]
  wire [11:0] idex_io_prev_csrAddr; // @[Core.scala 32:23]
  wire [31:0] idex_io_prev_csrData; // @[Core.scala 32:23]
  wire [3:0] idex_io_prev_excType; // @[Core.scala 32:23]
  wire [31:0] idex_io_prev_excValue; // @[Core.scala 32:23]
  wire  idex_io_prev_valid; // @[Core.scala 32:23]
  wire [31:0] idex_io_prev_inst; // @[Core.scala 32:23]
  wire [31:0] idex_io_prev_currentPc; // @[Core.scala 32:23]
  wire [3:0] idex_io_next_aluOp; // @[Core.scala 32:23]
  wire [31:0] idex_io_next_opr1; // @[Core.scala 32:23]
  wire [31:0] idex_io_next_opr2; // @[Core.scala 32:23]
  wire [3:0] idex_io_next_mduOp; // @[Core.scala 32:23]
  wire [4:0] idex_io_next_lsuOp; // @[Core.scala 32:23]
  wire [31:0] idex_io_next_lsuData; // @[Core.scala 32:23]
  wire  idex_io_next_regWen; // @[Core.scala 32:23]
  wire [4:0] idex_io_next_regWaddr; // @[Core.scala 32:23]
  wire [2:0] idex_io_next_csrOp; // @[Core.scala 32:23]
  wire [11:0] idex_io_next_csrAddr; // @[Core.scala 32:23]
  wire [31:0] idex_io_next_csrData; // @[Core.scala 32:23]
  wire [3:0] idex_io_next_excType; // @[Core.scala 32:23]
  wire [31:0] idex_io_next_excValue; // @[Core.scala 32:23]
  wire  idex_io_next_valid; // @[Core.scala 32:23]
  wire [31:0] idex_io_next_inst; // @[Core.scala 32:23]
  wire [31:0] idex_io_next_currentPc; // @[Core.scala 32:23]
  wire  alu_clock; // @[Core.scala 33:23]
  wire  alu_reset; // @[Core.scala 33:23]
  wire [3:0] alu_io_decoder_aluOp; // @[Core.scala 33:23]
  wire [31:0] alu_io_decoder_opr1; // @[Core.scala 33:23]
  wire [31:0] alu_io_decoder_opr2; // @[Core.scala 33:23]
  wire [3:0] alu_io_decoder_mduOp; // @[Core.scala 33:23]
  wire [4:0] alu_io_decoder_lsuOp; // @[Core.scala 33:23]
  wire [31:0] alu_io_decoder_lsuData; // @[Core.scala 33:23]
  wire  alu_io_decoder_regWen; // @[Core.scala 33:23]
  wire [4:0] alu_io_decoder_regWaddr; // @[Core.scala 33:23]
  wire [2:0] alu_io_decoder_csrOp; // @[Core.scala 33:23]
  wire [11:0] alu_io_decoder_csrAddr; // @[Core.scala 33:23]
  wire [31:0] alu_io_decoder_csrData; // @[Core.scala 33:23]
  wire [3:0] alu_io_decoder_excType; // @[Core.scala 33:23]
  wire [31:0] alu_io_decoder_excValue; // @[Core.scala 33:23]
  wire  alu_io_decoder_valid; // @[Core.scala 33:23]
  wire [31:0] alu_io_decoder_inst; // @[Core.scala 33:23]
  wire [31:0] alu_io_decoder_currentPc; // @[Core.scala 33:23]
  wire  alu_io_flush; // @[Core.scala 33:23]
  wire  alu_io_stallReq; // @[Core.scala 33:23]
  wire [2:0] alu_io_csrRead_op; // @[Core.scala 33:23]
  wire  alu_io_csrRead_valid; // @[Core.scala 33:23]
  wire [11:0] alu_io_csrRead_addr; // @[Core.scala 33:23]
  wire [31:0] alu_io_csrRead_data; // @[Core.scala 33:23]
  wire [4:0] alu_io_alu_lsuOp; // @[Core.scala 33:23]
  wire [31:0] alu_io_alu_lsuData; // @[Core.scala 33:23]
  wire  alu_io_alu_reg_en; // @[Core.scala 33:23]
  wire [4:0] alu_io_alu_reg_addr; // @[Core.scala 33:23]
  wire [31:0] alu_io_alu_reg_data; // @[Core.scala 33:23]
  wire  alu_io_alu_reg_load; // @[Core.scala 33:23]
  wire [2:0] alu_io_alu_csr_op; // @[Core.scala 33:23]
  wire [11:0] alu_io_alu_csr_addr; // @[Core.scala 33:23]
  wire [31:0] alu_io_alu_csr_data; // @[Core.scala 33:23]
  wire  alu_io_alu_csr_retired; // @[Core.scala 33:23]
  wire [3:0] alu_io_alu_excType; // @[Core.scala 33:23]
  wire [31:0] alu_io_alu_excValue; // @[Core.scala 33:23]
  wire  alu_io_alu_valid; // @[Core.scala 33:23]
  wire [31:0] alu_io_alu_inst; // @[Core.scala 33:23]
  wire [31:0] alu_io_alu_currentPc; // @[Core.scala 33:23]
  wire  exmem_clock; // @[Core.scala 34:23]
  wire  exmem_reset; // @[Core.scala 34:23]
  wire  exmem_io_flush; // @[Core.scala 34:23]
  wire  exmem_io_stallPrev; // @[Core.scala 34:23]
  wire  exmem_io_stallNext; // @[Core.scala 34:23]
  wire [4:0] exmem_io_prev_lsuOp; // @[Core.scala 34:23]
  wire [31:0] exmem_io_prev_lsuData; // @[Core.scala 34:23]
  wire  exmem_io_prev_reg_en; // @[Core.scala 34:23]
  wire [4:0] exmem_io_prev_reg_addr; // @[Core.scala 34:23]
  wire [31:0] exmem_io_prev_reg_data; // @[Core.scala 34:23]
  wire [2:0] exmem_io_prev_csr_op; // @[Core.scala 34:23]
  wire [11:0] exmem_io_prev_csr_addr; // @[Core.scala 34:23]
  wire [31:0] exmem_io_prev_csr_data; // @[Core.scala 34:23]
  wire  exmem_io_prev_csr_retired; // @[Core.scala 34:23]
  wire [3:0] exmem_io_prev_excType; // @[Core.scala 34:23]
  wire [31:0] exmem_io_prev_excValue; // @[Core.scala 34:23]
  wire  exmem_io_prev_valid; // @[Core.scala 34:23]
  wire [31:0] exmem_io_prev_inst; // @[Core.scala 34:23]
  wire [31:0] exmem_io_prev_currentPc; // @[Core.scala 34:23]
  wire [4:0] exmem_io_next_lsuOp; // @[Core.scala 34:23]
  wire [31:0] exmem_io_next_lsuData; // @[Core.scala 34:23]
  wire  exmem_io_next_reg_en; // @[Core.scala 34:23]
  wire [4:0] exmem_io_next_reg_addr; // @[Core.scala 34:23]
  wire [31:0] exmem_io_next_reg_data; // @[Core.scala 34:23]
  wire [2:0] exmem_io_next_csr_op; // @[Core.scala 34:23]
  wire [11:0] exmem_io_next_csr_addr; // @[Core.scala 34:23]
  wire [31:0] exmem_io_next_csr_data; // @[Core.scala 34:23]
  wire  exmem_io_next_csr_retired; // @[Core.scala 34:23]
  wire [3:0] exmem_io_next_excType; // @[Core.scala 34:23]
  wire [31:0] exmem_io_next_excValue; // @[Core.scala 34:23]
  wire  exmem_io_next_valid; // @[Core.scala 34:23]
  wire [31:0] exmem_io_next_inst; // @[Core.scala 34:23]
  wire [31:0] exmem_io_next_currentPc; // @[Core.scala 34:23]
  wire  mem_clock; // @[Core.scala 35:23]
  wire  mem_reset; // @[Core.scala 35:23]
  wire [4:0] mem_io_alu_lsuOp; // @[Core.scala 35:23]
  wire [31:0] mem_io_alu_lsuData; // @[Core.scala 35:23]
  wire  mem_io_alu_reg_en; // @[Core.scala 35:23]
  wire [4:0] mem_io_alu_reg_addr; // @[Core.scala 35:23]
  wire [31:0] mem_io_alu_reg_data; // @[Core.scala 35:23]
  wire [2:0] mem_io_alu_csr_op; // @[Core.scala 35:23]
  wire [11:0] mem_io_alu_csr_addr; // @[Core.scala 35:23]
  wire [31:0] mem_io_alu_csr_data; // @[Core.scala 35:23]
  wire  mem_io_alu_csr_retired; // @[Core.scala 35:23]
  wire [3:0] mem_io_alu_excType; // @[Core.scala 35:23]
  wire [31:0] mem_io_alu_excValue; // @[Core.scala 35:23]
  wire  mem_io_alu_valid; // @[Core.scala 35:23]
  wire [31:0] mem_io_alu_inst; // @[Core.scala 35:23]
  wire [31:0] mem_io_alu_currentPc; // @[Core.scala 35:23]
  wire  mem_io_flush; // @[Core.scala 35:23]
  wire  mem_io_stallReq; // @[Core.scala 35:23]
  wire  mem_io_flushReq; // @[Core.scala 35:23]
  wire [31:0] mem_io_flushPc; // @[Core.scala 35:23]
  wire  mem_io_ram_en; // @[Core.scala 35:23]
  wire  mem_io_ram_valid; // @[Core.scala 35:23]
  wire  mem_io_ram_fault; // @[Core.scala 35:23]
  wire [3:0] mem_io_ram_wen; // @[Core.scala 35:23]
  wire [31:0] mem_io_ram_addr; // @[Core.scala 35:23]
  wire [31:0] mem_io_ram_rdata; // @[Core.scala 35:23]
  wire [31:0] mem_io_ram_wdata; // @[Core.scala 35:23]
  wire  mem_io_flushIc; // @[Core.scala 35:23]
  wire  mem_io_flushDc; // @[Core.scala 35:23]
  wire  mem_io_flushIt; // @[Core.scala 35:23]
  wire  mem_io_flushDt; // @[Core.scala 35:23]
  wire  mem_io_csrHasInt; // @[Core.scala 35:23]
  wire  mem_io_csrBusy; // @[Core.scala 35:23]
  wire [1:0] mem_io_csrMode; // @[Core.scala 35:23]
  wire [31:0] mem_io_excMon_addr; // @[Core.scala 35:23]
  wire  mem_io_excMon_valid; // @[Core.scala 35:23]
  wire  mem_io_except_hasTrap; // @[Core.scala 35:23]
  wire  mem_io_except_isSret; // @[Core.scala 35:23]
  wire  mem_io_except_isMret; // @[Core.scala 35:23]
  wire [30:0] mem_io_except_excCause; // @[Core.scala 35:23]
  wire [31:0] mem_io_except_excPc; // @[Core.scala 35:23]
  wire [31:0] mem_io_except_excValue; // @[Core.scala 35:23]
  wire  mem_io_mem_reg_en; // @[Core.scala 35:23]
  wire [4:0] mem_io_mem_reg_addr; // @[Core.scala 35:23]
  wire [31:0] mem_io_mem_reg_data; // @[Core.scala 35:23]
  wire  mem_io_mem_reg_load; // @[Core.scala 35:23]
  wire  mem_io_mem_memSigned; // @[Core.scala 35:23]
  wire [1:0] mem_io_mem_memSel; // @[Core.scala 35:23]
  wire [1:0] mem_io_mem_memWidth; // @[Core.scala 35:23]
  wire [2:0] mem_io_mem_csr_op; // @[Core.scala 35:23]
  wire [11:0] mem_io_mem_csr_addr; // @[Core.scala 35:23]
  wire [31:0] mem_io_mem_csr_data; // @[Core.scala 35:23]
  wire  mem_io_mem_csr_retired; // @[Core.scala 35:23]
  wire [31:0] mem_io_mem_excMon_addr; // @[Core.scala 35:23]
  wire  mem_io_mem_excMon_set; // @[Core.scala 35:23]
  wire  mem_io_mem_excMon_clear; // @[Core.scala 35:23]
  wire [31:0] mem_io_mem_currentPc; // @[Core.scala 35:23]
  wire  memwb_clock; // @[Core.scala 36:23]
  wire  memwb_reset; // @[Core.scala 36:23]
  wire  memwb_io_flush; // @[Core.scala 36:23]
  wire  memwb_io_stallPrev; // @[Core.scala 36:23]
  wire  memwb_io_stallNext; // @[Core.scala 36:23]
  wire  memwb_io_prev_reg_en; // @[Core.scala 36:23]
  wire [4:0] memwb_io_prev_reg_addr; // @[Core.scala 36:23]
  wire [31:0] memwb_io_prev_reg_data; // @[Core.scala 36:23]
  wire  memwb_io_prev_reg_load; // @[Core.scala 36:23]
  wire  memwb_io_prev_memSigned; // @[Core.scala 36:23]
  wire [1:0] memwb_io_prev_memSel; // @[Core.scala 36:23]
  wire [1:0] memwb_io_prev_memWidth; // @[Core.scala 36:23]
  wire [2:0] memwb_io_prev_csr_op; // @[Core.scala 36:23]
  wire [11:0] memwb_io_prev_csr_addr; // @[Core.scala 36:23]
  wire [31:0] memwb_io_prev_csr_data; // @[Core.scala 36:23]
  wire  memwb_io_prev_csr_retired; // @[Core.scala 36:23]
  wire [31:0] memwb_io_prev_excMon_addr; // @[Core.scala 36:23]
  wire  memwb_io_prev_excMon_set; // @[Core.scala 36:23]
  wire  memwb_io_prev_excMon_clear; // @[Core.scala 36:23]
  wire [31:0] memwb_io_prev_currentPc; // @[Core.scala 36:23]
  wire  memwb_io_next_reg_en; // @[Core.scala 36:23]
  wire [4:0] memwb_io_next_reg_addr; // @[Core.scala 36:23]
  wire [31:0] memwb_io_next_reg_data; // @[Core.scala 36:23]
  wire  memwb_io_next_reg_load; // @[Core.scala 36:23]
  wire  memwb_io_next_memSigned; // @[Core.scala 36:23]
  wire [1:0] memwb_io_next_memSel; // @[Core.scala 36:23]
  wire [1:0] memwb_io_next_memWidth; // @[Core.scala 36:23]
  wire [2:0] memwb_io_next_csr_op; // @[Core.scala 36:23]
  wire [11:0] memwb_io_next_csr_addr; // @[Core.scala 36:23]
  wire [31:0] memwb_io_next_csr_data; // @[Core.scala 36:23]
  wire  memwb_io_next_csr_retired; // @[Core.scala 36:23]
  wire [31:0] memwb_io_next_excMon_addr; // @[Core.scala 36:23]
  wire  memwb_io_next_excMon_set; // @[Core.scala 36:23]
  wire  memwb_io_next_excMon_clear; // @[Core.scala 36:23]
  wire [31:0] memwb_io_next_currentPc; // @[Core.scala 36:23]
  wire  wb_io_mem_reg_en; // @[Core.scala 37:23]
  wire [4:0] wb_io_mem_reg_addr; // @[Core.scala 37:23]
  wire [31:0] wb_io_mem_reg_data; // @[Core.scala 37:23]
  wire  wb_io_mem_reg_load; // @[Core.scala 37:23]
  wire  wb_io_mem_memSigned; // @[Core.scala 37:23]
  wire [1:0] wb_io_mem_memSel; // @[Core.scala 37:23]
  wire [1:0] wb_io_mem_memWidth; // @[Core.scala 37:23]
  wire [2:0] wb_io_mem_csr_op; // @[Core.scala 37:23]
  wire [11:0] wb_io_mem_csr_addr; // @[Core.scala 37:23]
  wire [31:0] wb_io_mem_csr_data; // @[Core.scala 37:23]
  wire  wb_io_mem_csr_retired; // @[Core.scala 37:23]
  wire [31:0] wb_io_mem_excMon_addr; // @[Core.scala 37:23]
  wire  wb_io_mem_excMon_set; // @[Core.scala 37:23]
  wire  wb_io_mem_excMon_clear; // @[Core.scala 37:23]
  wire [31:0] wb_io_mem_currentPc; // @[Core.scala 37:23]
  wire [31:0] wb_io_ramData; // @[Core.scala 37:23]
  wire  wb_io_reg_en; // @[Core.scala 37:23]
  wire [4:0] wb_io_reg_addr; // @[Core.scala 37:23]
  wire [31:0] wb_io_reg_data; // @[Core.scala 37:23]
  wire [2:0] wb_io_csr_op; // @[Core.scala 37:23]
  wire [11:0] wb_io_csr_addr; // @[Core.scala 37:23]
  wire [31:0] wb_io_csr_data; // @[Core.scala 37:23]
  wire  wb_io_csr_retired; // @[Core.scala 37:23]
  wire [31:0] wb_io_excMon_addr; // @[Core.scala 37:23]
  wire  wb_io_excMon_set; // @[Core.scala 37:23]
  wire  wb_io_excMon_clear; // @[Core.scala 37:23]
  wire  wb_io_debug_regWen; // @[Core.scala 37:23]
  wire [4:0] wb_io_debug_regWaddr; // @[Core.scala 37:23]
  wire [31:0] wb_io_debug_regWdata; // @[Core.scala 37:23]
  wire [31:0] wb_io_debug_pc; // @[Core.scala 37:23]
  wire  regfile_clock; // @[Core.scala 40:23]
  wire  regfile_reset; // @[Core.scala 40:23]
  wire  regfile_io_read1_en; // @[Core.scala 40:23]
  wire [4:0] regfile_io_read1_addr; // @[Core.scala 40:23]
  wire [31:0] regfile_io_read1_data; // @[Core.scala 40:23]
  wire  regfile_io_read2_en; // @[Core.scala 40:23]
  wire [4:0] regfile_io_read2_addr; // @[Core.scala 40:23]
  wire [31:0] regfile_io_read2_data; // @[Core.scala 40:23]
  wire  regfile_io_write_en; // @[Core.scala 40:23]
  wire [4:0] regfile_io_write_addr; // @[Core.scala 40:23]
  wire [31:0] regfile_io_write_data; // @[Core.scala 40:23]
  wire  csrfile_clock; // @[Core.scala 43:23]
  wire  csrfile_reset; // @[Core.scala 43:23]
  wire [2:0] csrfile_io_read_op; // @[Core.scala 43:23]
  wire  csrfile_io_read_valid; // @[Core.scala 43:23]
  wire [11:0] csrfile_io_read_addr; // @[Core.scala 43:23]
  wire [31:0] csrfile_io_read_data; // @[Core.scala 43:23]
  wire [2:0] csrfile_io_write_op; // @[Core.scala 43:23]
  wire [11:0] csrfile_io_write_addr; // @[Core.scala 43:23]
  wire [31:0] csrfile_io_write_data; // @[Core.scala 43:23]
  wire  csrfile_io_write_retired; // @[Core.scala 43:23]
  wire  csrfile_io_irq_timer; // @[Core.scala 43:23]
  wire  csrfile_io_irq_soft; // @[Core.scala 43:23]
  wire  csrfile_io_irq_extern; // @[Core.scala 43:23]
  wire  csrfile_io_except_hasTrap; // @[Core.scala 43:23]
  wire  csrfile_io_except_isSret; // @[Core.scala 43:23]
  wire  csrfile_io_except_isMret; // @[Core.scala 43:23]
  wire [30:0] csrfile_io_except_excCause; // @[Core.scala 43:23]
  wire [31:0] csrfile_io_except_excPc; // @[Core.scala 43:23]
  wire [31:0] csrfile_io_except_excValue; // @[Core.scala 43:23]
  wire  csrfile_io_hasInt; // @[Core.scala 43:23]
  wire  csrfile_io_busy; // @[Core.scala 43:23]
  wire [1:0] csrfile_io_mode; // @[Core.scala 43:23]
  wire [31:0] csrfile_io_sepc; // @[Core.scala 43:23]
  wire [31:0] csrfile_io_mepc; // @[Core.scala 43:23]
  wire [31:0] csrfile_io_trapVec; // @[Core.scala 43:23]
  wire  csrfile_io_pageEn; // @[Core.scala 43:23]
  wire [21:0] csrfile_io_basePpn; // @[Core.scala 43:23]
  wire  csrfile_io_sum; // @[Core.scala 43:23]
  wire  excMon_clock; // @[Core.scala 46:23]
  wire  excMon_reset; // @[Core.scala 46:23]
  wire  excMon_io_flush; // @[Core.scala 46:23]
  wire [31:0] excMon_io_check_addr; // @[Core.scala 46:23]
  wire  excMon_io_check_valid; // @[Core.scala 46:23]
  wire [31:0] excMon_io_update_addr; // @[Core.scala 46:23]
  wire  excMon_io_update_set; // @[Core.scala 46:23]
  wire  excMon_io_update_clear; // @[Core.scala 46:23]
  wire  resolve_io_regRead1_en; // @[Core.scala 49:23]
  wire [4:0] resolve_io_regRead1_addr; // @[Core.scala 49:23]
  wire [31:0] resolve_io_regRead1_data; // @[Core.scala 49:23]
  wire  resolve_io_regRead2_en; // @[Core.scala 49:23]
  wire [4:0] resolve_io_regRead2_addr; // @[Core.scala 49:23]
  wire [31:0] resolve_io_regRead2_data; // @[Core.scala 49:23]
  wire [2:0] resolve_io_csrRead_op; // @[Core.scala 49:23]
  wire  resolve_io_csrRead_valid; // @[Core.scala 49:23]
  wire [11:0] resolve_io_csrRead_addr; // @[Core.scala 49:23]
  wire [31:0] resolve_io_csrRead_data; // @[Core.scala 49:23]
  wire [31:0] resolve_io_check_addr; // @[Core.scala 49:23]
  wire  resolve_io_check_valid; // @[Core.scala 49:23]
  wire  resolve_io_aluReg_en; // @[Core.scala 49:23]
  wire [4:0] resolve_io_aluReg_addr; // @[Core.scala 49:23]
  wire [31:0] resolve_io_aluReg_data; // @[Core.scala 49:23]
  wire  resolve_io_aluReg_load; // @[Core.scala 49:23]
  wire  resolve_io_memReg_en; // @[Core.scala 49:23]
  wire [4:0] resolve_io_memReg_addr; // @[Core.scala 49:23]
  wire [31:0] resolve_io_memReg_data; // @[Core.scala 49:23]
  wire  resolve_io_memReg_load; // @[Core.scala 49:23]
  wire [2:0] resolve_io_memCsr_op; // @[Core.scala 49:23]
  wire [11:0] resolve_io_memCsr_addr; // @[Core.scala 49:23]
  wire  resolve_io_wbReg_en; // @[Core.scala 49:23]
  wire [4:0] resolve_io_wbReg_addr; // @[Core.scala 49:23]
  wire [31:0] resolve_io_wbReg_data; // @[Core.scala 49:23]
  wire [2:0] resolve_io_wbCsr_op; // @[Core.scala 49:23]
  wire [11:0] resolve_io_wbCsr_addr; // @[Core.scala 49:23]
  wire [31:0] resolve_io_wbExcMon_addr; // @[Core.scala 49:23]
  wire  resolve_io_wbExcMon_set; // @[Core.scala 49:23]
  wire  resolve_io_wbExcMon_clear; // @[Core.scala 49:23]
  wire  resolve_io_rf1_en; // @[Core.scala 49:23]
  wire [4:0] resolve_io_rf1_addr; // @[Core.scala 49:23]
  wire [31:0] resolve_io_rf1_data; // @[Core.scala 49:23]
  wire  resolve_io_rf2_en; // @[Core.scala 49:23]
  wire [4:0] resolve_io_rf2_addr; // @[Core.scala 49:23]
  wire [31:0] resolve_io_rf2_data; // @[Core.scala 49:23]
  wire [2:0] resolve_io_csr_op; // @[Core.scala 49:23]
  wire  resolve_io_csr_valid; // @[Core.scala 49:23]
  wire [11:0] resolve_io_csr_addr; // @[Core.scala 49:23]
  wire [31:0] resolve_io_csr_data; // @[Core.scala 49:23]
  wire [31:0] resolve_io_excMon_addr; // @[Core.scala 49:23]
  wire  resolve_io_excMon_valid; // @[Core.scala 49:23]
  wire  resolve_io_loadFlag; // @[Core.scala 49:23]
  wire  resolve_io_csrFlag; // @[Core.scala 49:23]
  wire  control_io_fetch; // @[Core.scala 50:23]
  wire  control_io_alu; // @[Core.scala 50:23]
  wire  control_io_mem; // @[Core.scala 50:23]
  wire  control_io_decFlush; // @[Core.scala 50:23]
  wire [31:0] control_io_decTarget; // @[Core.scala 50:23]
  wire  control_io_memFlush; // @[Core.scala 50:23]
  wire [31:0] control_io_memTarget; // @[Core.scala 50:23]
  wire  control_io_load; // @[Core.scala 50:23]
  wire  control_io_csr; // @[Core.scala 50:23]
  wire  control_io_except_hasTrap; // @[Core.scala 50:23]
  wire  control_io_except_isSret; // @[Core.scala 50:23]
  wire  control_io_except_isMret; // @[Core.scala 50:23]
  wire [31:0] control_io_csrSepc; // @[Core.scala 50:23]
  wire [31:0] control_io_csrMepc; // @[Core.scala 50:23]
  wire [31:0] control_io_csrTvec; // @[Core.scala 50:23]
  wire  control_io_stallIf; // @[Core.scala 50:23]
  wire  control_io_stallId; // @[Core.scala 50:23]
  wire  control_io_stallEx; // @[Core.scala 50:23]
  wire  control_io_stallMm; // @[Core.scala 50:23]
  wire  control_io_stallWb; // @[Core.scala 50:23]
  wire  control_io_flush; // @[Core.scala 50:23]
  wire  control_io_flushIf; // @[Core.scala 50:23]
  wire [31:0] control_io_flushPc; // @[Core.scala 50:23]
  Fetch fetch ( // @[Core.scala 29:23]
    .clock(fetch_clock),
    .reset(fetch_reset),
    .io_flush(fetch_io_flush),
    .io_stall(fetch_io_stall),
    .io_stallReq(fetch_io_stallReq),
    .io_flushPc(fetch_io_flushPc),
    .io_rom_valid(fetch_io_rom_valid),
    .io_rom_fault(fetch_io_rom_fault),
    .io_rom_addr(fetch_io_rom_addr),
    .io_branch_branch(fetch_io_branch_branch),
    .io_branch_jump(fetch_io_branch_jump),
    .io_branch_taken(fetch_io_branch_taken),
    .io_branch_index(fetch_io_branch_index),
    .io_branch_pc(fetch_io_branch_pc),
    .io_branch_target(fetch_io_branch_target),
    .io_fetch_valid(fetch_io_fetch_valid),
    .io_fetch_pc(fetch_io_fetch_pc),
    .io_fetch_taken(fetch_io_fetch_taken),
    .io_fetch_target(fetch_io_fetch_target),
    .io_fetch_predIndex(fetch_io_fetch_predIndex),
    .io_fetch_pageFault(fetch_io_fetch_pageFault)
  );
  MidStage ifid ( // @[Core.scala 30:23]
    .clock(ifid_clock),
    .reset(ifid_reset),
    .io_flush(ifid_io_flush),
    .io_stallPrev(ifid_io_stallPrev),
    .io_stallNext(ifid_io_stallNext),
    .io_prev_valid(ifid_io_prev_valid),
    .io_prev_pc(ifid_io_prev_pc),
    .io_prev_taken(ifid_io_prev_taken),
    .io_prev_target(ifid_io_prev_target),
    .io_prev_predIndex(ifid_io_prev_predIndex),
    .io_prev_pageFault(ifid_io_prev_pageFault),
    .io_next_valid(ifid_io_next_valid),
    .io_next_pc(ifid_io_next_pc),
    .io_next_taken(ifid_io_next_taken),
    .io_next_target(ifid_io_next_target),
    .io_next_predIndex(ifid_io_next_predIndex),
    .io_next_pageFault(ifid_io_next_pageFault)
  );
  Decoder decoder ( // @[Core.scala 31:23]
    .clock(decoder_clock),
    .io_fetch_valid(decoder_io_fetch_valid),
    .io_fetch_pc(decoder_io_fetch_pc),
    .io_fetch_taken(decoder_io_fetch_taken),
    .io_fetch_target(decoder_io_fetch_target),
    .io_fetch_predIndex(decoder_io_fetch_predIndex),
    .io_fetch_pageFault(decoder_io_fetch_pageFault),
    .io_inst(decoder_io_inst),
    .io_stallId(decoder_io_stallId),
    .io_flushIf(decoder_io_flushIf),
    .io_flushPc(decoder_io_flushPc),
    .io_read1_en(decoder_io_read1_en),
    .io_read1_addr(decoder_io_read1_addr),
    .io_read1_data(decoder_io_read1_data),
    .io_read2_en(decoder_io_read2_en),
    .io_read2_addr(decoder_io_read2_addr),
    .io_read2_data(decoder_io_read2_data),
    .io_branch_branch(decoder_io_branch_branch),
    .io_branch_jump(decoder_io_branch_jump),
    .io_branch_taken(decoder_io_branch_taken),
    .io_branch_index(decoder_io_branch_index),
    .io_branch_pc(decoder_io_branch_pc),
    .io_branch_target(decoder_io_branch_target),
    .io_decoder_aluOp(decoder_io_decoder_aluOp),
    .io_decoder_opr1(decoder_io_decoder_opr1),
    .io_decoder_opr2(decoder_io_decoder_opr2),
    .io_decoder_mduOp(decoder_io_decoder_mduOp),
    .io_decoder_lsuOp(decoder_io_decoder_lsuOp),
    .io_decoder_lsuData(decoder_io_decoder_lsuData),
    .io_decoder_regWen(decoder_io_decoder_regWen),
    .io_decoder_regWaddr(decoder_io_decoder_regWaddr),
    .io_decoder_csrOp(decoder_io_decoder_csrOp),
    .io_decoder_csrAddr(decoder_io_decoder_csrAddr),
    .io_decoder_csrData(decoder_io_decoder_csrData),
    .io_decoder_excType(decoder_io_decoder_excType),
    .io_decoder_excValue(decoder_io_decoder_excValue),
    .io_decoder_valid(decoder_io_decoder_valid),
    .io_decoder_inst(decoder_io_decoder_inst),
    .io_decoder_currentPc(decoder_io_decoder_currentPc)
  );
  MidStage_1 idex ( // @[Core.scala 32:23]
    .clock(idex_clock),
    .reset(idex_reset),
    .io_flush(idex_io_flush),
    .io_stallPrev(idex_io_stallPrev),
    .io_stallNext(idex_io_stallNext),
    .io_prev_aluOp(idex_io_prev_aluOp),
    .io_prev_opr1(idex_io_prev_opr1),
    .io_prev_opr2(idex_io_prev_opr2),
    .io_prev_mduOp(idex_io_prev_mduOp),
    .io_prev_lsuOp(idex_io_prev_lsuOp),
    .io_prev_lsuData(idex_io_prev_lsuData),
    .io_prev_regWen(idex_io_prev_regWen),
    .io_prev_regWaddr(idex_io_prev_regWaddr),
    .io_prev_csrOp(idex_io_prev_csrOp),
    .io_prev_csrAddr(idex_io_prev_csrAddr),
    .io_prev_csrData(idex_io_prev_csrData),
    .io_prev_excType(idex_io_prev_excType),
    .io_prev_excValue(idex_io_prev_excValue),
    .io_prev_valid(idex_io_prev_valid),
    .io_prev_inst(idex_io_prev_inst),
    .io_prev_currentPc(idex_io_prev_currentPc),
    .io_next_aluOp(idex_io_next_aluOp),
    .io_next_opr1(idex_io_next_opr1),
    .io_next_opr2(idex_io_next_opr2),
    .io_next_mduOp(idex_io_next_mduOp),
    .io_next_lsuOp(idex_io_next_lsuOp),
    .io_next_lsuData(idex_io_next_lsuData),
    .io_next_regWen(idex_io_next_regWen),
    .io_next_regWaddr(idex_io_next_regWaddr),
    .io_next_csrOp(idex_io_next_csrOp),
    .io_next_csrAddr(idex_io_next_csrAddr),
    .io_next_csrData(idex_io_next_csrData),
    .io_next_excType(idex_io_next_excType),
    .io_next_excValue(idex_io_next_excValue),
    .io_next_valid(idex_io_next_valid),
    .io_next_inst(idex_io_next_inst),
    .io_next_currentPc(idex_io_next_currentPc)
  );
  ALU alu ( // @[Core.scala 33:23]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_decoder_aluOp(alu_io_decoder_aluOp),
    .io_decoder_opr1(alu_io_decoder_opr1),
    .io_decoder_opr2(alu_io_decoder_opr2),
    .io_decoder_mduOp(alu_io_decoder_mduOp),
    .io_decoder_lsuOp(alu_io_decoder_lsuOp),
    .io_decoder_lsuData(alu_io_decoder_lsuData),
    .io_decoder_regWen(alu_io_decoder_regWen),
    .io_decoder_regWaddr(alu_io_decoder_regWaddr),
    .io_decoder_csrOp(alu_io_decoder_csrOp),
    .io_decoder_csrAddr(alu_io_decoder_csrAddr),
    .io_decoder_csrData(alu_io_decoder_csrData),
    .io_decoder_excType(alu_io_decoder_excType),
    .io_decoder_excValue(alu_io_decoder_excValue),
    .io_decoder_valid(alu_io_decoder_valid),
    .io_decoder_inst(alu_io_decoder_inst),
    .io_decoder_currentPc(alu_io_decoder_currentPc),
    .io_flush(alu_io_flush),
    .io_stallReq(alu_io_stallReq),
    .io_csrRead_op(alu_io_csrRead_op),
    .io_csrRead_valid(alu_io_csrRead_valid),
    .io_csrRead_addr(alu_io_csrRead_addr),
    .io_csrRead_data(alu_io_csrRead_data),
    .io_alu_lsuOp(alu_io_alu_lsuOp),
    .io_alu_lsuData(alu_io_alu_lsuData),
    .io_alu_reg_en(alu_io_alu_reg_en),
    .io_alu_reg_addr(alu_io_alu_reg_addr),
    .io_alu_reg_data(alu_io_alu_reg_data),
    .io_alu_reg_load(alu_io_alu_reg_load),
    .io_alu_csr_op(alu_io_alu_csr_op),
    .io_alu_csr_addr(alu_io_alu_csr_addr),
    .io_alu_csr_data(alu_io_alu_csr_data),
    .io_alu_csr_retired(alu_io_alu_csr_retired),
    .io_alu_excType(alu_io_alu_excType),
    .io_alu_excValue(alu_io_alu_excValue),
    .io_alu_valid(alu_io_alu_valid),
    .io_alu_inst(alu_io_alu_inst),
    .io_alu_currentPc(alu_io_alu_currentPc)
  );
  MidStage_2 exmem ( // @[Core.scala 34:23]
    .clock(exmem_clock),
    .reset(exmem_reset),
    .io_flush(exmem_io_flush),
    .io_stallPrev(exmem_io_stallPrev),
    .io_stallNext(exmem_io_stallNext),
    .io_prev_lsuOp(exmem_io_prev_lsuOp),
    .io_prev_lsuData(exmem_io_prev_lsuData),
    .io_prev_reg_en(exmem_io_prev_reg_en),
    .io_prev_reg_addr(exmem_io_prev_reg_addr),
    .io_prev_reg_data(exmem_io_prev_reg_data),
    .io_prev_csr_op(exmem_io_prev_csr_op),
    .io_prev_csr_addr(exmem_io_prev_csr_addr),
    .io_prev_csr_data(exmem_io_prev_csr_data),
    .io_prev_csr_retired(exmem_io_prev_csr_retired),
    .io_prev_excType(exmem_io_prev_excType),
    .io_prev_excValue(exmem_io_prev_excValue),
    .io_prev_valid(exmem_io_prev_valid),
    .io_prev_inst(exmem_io_prev_inst),
    .io_prev_currentPc(exmem_io_prev_currentPc),
    .io_next_lsuOp(exmem_io_next_lsuOp),
    .io_next_lsuData(exmem_io_next_lsuData),
    .io_next_reg_en(exmem_io_next_reg_en),
    .io_next_reg_addr(exmem_io_next_reg_addr),
    .io_next_reg_data(exmem_io_next_reg_data),
    .io_next_csr_op(exmem_io_next_csr_op),
    .io_next_csr_addr(exmem_io_next_csr_addr),
    .io_next_csr_data(exmem_io_next_csr_data),
    .io_next_csr_retired(exmem_io_next_csr_retired),
    .io_next_excType(exmem_io_next_excType),
    .io_next_excValue(exmem_io_next_excValue),
    .io_next_valid(exmem_io_next_valid),
    .io_next_inst(exmem_io_next_inst),
    .io_next_currentPc(exmem_io_next_currentPc)
  );
  Mem mem ( // @[Core.scala 35:23]
    .clock(mem_clock),
    .reset(mem_reset),
    .io_alu_lsuOp(mem_io_alu_lsuOp),
    .io_alu_lsuData(mem_io_alu_lsuData),
    .io_alu_reg_en(mem_io_alu_reg_en),
    .io_alu_reg_addr(mem_io_alu_reg_addr),
    .io_alu_reg_data(mem_io_alu_reg_data),
    .io_alu_csr_op(mem_io_alu_csr_op),
    .io_alu_csr_addr(mem_io_alu_csr_addr),
    .io_alu_csr_data(mem_io_alu_csr_data),
    .io_alu_csr_retired(mem_io_alu_csr_retired),
    .io_alu_excType(mem_io_alu_excType),
    .io_alu_excValue(mem_io_alu_excValue),
    .io_alu_valid(mem_io_alu_valid),
    .io_alu_inst(mem_io_alu_inst),
    .io_alu_currentPc(mem_io_alu_currentPc),
    .io_flush(mem_io_flush),
    .io_stallReq(mem_io_stallReq),
    .io_flushReq(mem_io_flushReq),
    .io_flushPc(mem_io_flushPc),
    .io_ram_en(mem_io_ram_en),
    .io_ram_valid(mem_io_ram_valid),
    .io_ram_fault(mem_io_ram_fault),
    .io_ram_wen(mem_io_ram_wen),
    .io_ram_addr(mem_io_ram_addr),
    .io_ram_rdata(mem_io_ram_rdata),
    .io_ram_wdata(mem_io_ram_wdata),
    .io_flushIc(mem_io_flushIc),
    .io_flushDc(mem_io_flushDc),
    .io_flushIt(mem_io_flushIt),
    .io_flushDt(mem_io_flushDt),
    .io_csrHasInt(mem_io_csrHasInt),
    .io_csrBusy(mem_io_csrBusy),
    .io_csrMode(mem_io_csrMode),
    .io_excMon_addr(mem_io_excMon_addr),
    .io_excMon_valid(mem_io_excMon_valid),
    .io_except_hasTrap(mem_io_except_hasTrap),
    .io_except_isSret(mem_io_except_isSret),
    .io_except_isMret(mem_io_except_isMret),
    .io_except_excCause(mem_io_except_excCause),
    .io_except_excPc(mem_io_except_excPc),
    .io_except_excValue(mem_io_except_excValue),
    .io_mem_reg_en(mem_io_mem_reg_en),
    .io_mem_reg_addr(mem_io_mem_reg_addr),
    .io_mem_reg_data(mem_io_mem_reg_data),
    .io_mem_reg_load(mem_io_mem_reg_load),
    .io_mem_memSigned(mem_io_mem_memSigned),
    .io_mem_memSel(mem_io_mem_memSel),
    .io_mem_memWidth(mem_io_mem_memWidth),
    .io_mem_csr_op(mem_io_mem_csr_op),
    .io_mem_csr_addr(mem_io_mem_csr_addr),
    .io_mem_csr_data(mem_io_mem_csr_data),
    .io_mem_csr_retired(mem_io_mem_csr_retired),
    .io_mem_excMon_addr(mem_io_mem_excMon_addr),
    .io_mem_excMon_set(mem_io_mem_excMon_set),
    .io_mem_excMon_clear(mem_io_mem_excMon_clear),
    .io_mem_currentPc(mem_io_mem_currentPc)
  );
  MidStage_3 memwb ( // @[Core.scala 36:23]
    .clock(memwb_clock),
    .reset(memwb_reset),
    .io_flush(memwb_io_flush),
    .io_stallPrev(memwb_io_stallPrev),
    .io_stallNext(memwb_io_stallNext),
    .io_prev_reg_en(memwb_io_prev_reg_en),
    .io_prev_reg_addr(memwb_io_prev_reg_addr),
    .io_prev_reg_data(memwb_io_prev_reg_data),
    .io_prev_reg_load(memwb_io_prev_reg_load),
    .io_prev_memSigned(memwb_io_prev_memSigned),
    .io_prev_memSel(memwb_io_prev_memSel),
    .io_prev_memWidth(memwb_io_prev_memWidth),
    .io_prev_csr_op(memwb_io_prev_csr_op),
    .io_prev_csr_addr(memwb_io_prev_csr_addr),
    .io_prev_csr_data(memwb_io_prev_csr_data),
    .io_prev_csr_retired(memwb_io_prev_csr_retired),
    .io_prev_excMon_addr(memwb_io_prev_excMon_addr),
    .io_prev_excMon_set(memwb_io_prev_excMon_set),
    .io_prev_excMon_clear(memwb_io_prev_excMon_clear),
    .io_prev_currentPc(memwb_io_prev_currentPc),
    .io_next_reg_en(memwb_io_next_reg_en),
    .io_next_reg_addr(memwb_io_next_reg_addr),
    .io_next_reg_data(memwb_io_next_reg_data),
    .io_next_reg_load(memwb_io_next_reg_load),
    .io_next_memSigned(memwb_io_next_memSigned),
    .io_next_memSel(memwb_io_next_memSel),
    .io_next_memWidth(memwb_io_next_memWidth),
    .io_next_csr_op(memwb_io_next_csr_op),
    .io_next_csr_addr(memwb_io_next_csr_addr),
    .io_next_csr_data(memwb_io_next_csr_data),
    .io_next_csr_retired(memwb_io_next_csr_retired),
    .io_next_excMon_addr(memwb_io_next_excMon_addr),
    .io_next_excMon_set(memwb_io_next_excMon_set),
    .io_next_excMon_clear(memwb_io_next_excMon_clear),
    .io_next_currentPc(memwb_io_next_currentPc)
  );
  WriteBack wb ( // @[Core.scala 37:23]
    .io_mem_reg_en(wb_io_mem_reg_en),
    .io_mem_reg_addr(wb_io_mem_reg_addr),
    .io_mem_reg_data(wb_io_mem_reg_data),
    .io_mem_reg_load(wb_io_mem_reg_load),
    .io_mem_memSigned(wb_io_mem_memSigned),
    .io_mem_memSel(wb_io_mem_memSel),
    .io_mem_memWidth(wb_io_mem_memWidth),
    .io_mem_csr_op(wb_io_mem_csr_op),
    .io_mem_csr_addr(wb_io_mem_csr_addr),
    .io_mem_csr_data(wb_io_mem_csr_data),
    .io_mem_csr_retired(wb_io_mem_csr_retired),
    .io_mem_excMon_addr(wb_io_mem_excMon_addr),
    .io_mem_excMon_set(wb_io_mem_excMon_set),
    .io_mem_excMon_clear(wb_io_mem_excMon_clear),
    .io_mem_currentPc(wb_io_mem_currentPc),
    .io_ramData(wb_io_ramData),
    .io_reg_en(wb_io_reg_en),
    .io_reg_addr(wb_io_reg_addr),
    .io_reg_data(wb_io_reg_data),
    .io_csr_op(wb_io_csr_op),
    .io_csr_addr(wb_io_csr_addr),
    .io_csr_data(wb_io_csr_data),
    .io_csr_retired(wb_io_csr_retired),
    .io_excMon_addr(wb_io_excMon_addr),
    .io_excMon_set(wb_io_excMon_set),
    .io_excMon_clear(wb_io_excMon_clear),
    .io_debug_regWen(wb_io_debug_regWen),
    .io_debug_regWaddr(wb_io_debug_regWaddr),
    .io_debug_regWdata(wb_io_debug_regWdata),
    .io_debug_pc(wb_io_debug_pc)
  );
  RegFile regfile ( // @[Core.scala 40:23]
    .clock(regfile_clock),
    .reset(regfile_reset),
    .io_read1_en(regfile_io_read1_en),
    .io_read1_addr(regfile_io_read1_addr),
    .io_read1_data(regfile_io_read1_data),
    .io_read2_en(regfile_io_read2_en),
    .io_read2_addr(regfile_io_read2_addr),
    .io_read2_data(regfile_io_read2_data),
    .io_write_en(regfile_io_write_en),
    .io_write_addr(regfile_io_write_addr),
    .io_write_data(regfile_io_write_data)
  );
  CsrFile csrfile ( // @[Core.scala 43:23]
    .clock(csrfile_clock),
    .reset(csrfile_reset),
    .io_read_op(csrfile_io_read_op),
    .io_read_valid(csrfile_io_read_valid),
    .io_read_addr(csrfile_io_read_addr),
    .io_read_data(csrfile_io_read_data),
    .io_write_op(csrfile_io_write_op),
    .io_write_addr(csrfile_io_write_addr),
    .io_write_data(csrfile_io_write_data),
    .io_write_retired(csrfile_io_write_retired),
    .io_irq_timer(csrfile_io_irq_timer),
    .io_irq_soft(csrfile_io_irq_soft),
    .io_irq_extern(csrfile_io_irq_extern),
    .io_except_hasTrap(csrfile_io_except_hasTrap),
    .io_except_isSret(csrfile_io_except_isSret),
    .io_except_isMret(csrfile_io_except_isMret),
    .io_except_excCause(csrfile_io_except_excCause),
    .io_except_excPc(csrfile_io_except_excPc),
    .io_except_excValue(csrfile_io_except_excValue),
    .io_hasInt(csrfile_io_hasInt),
    .io_busy(csrfile_io_busy),
    .io_mode(csrfile_io_mode),
    .io_sepc(csrfile_io_sepc),
    .io_mepc(csrfile_io_mepc),
    .io_trapVec(csrfile_io_trapVec),
    .io_pageEn(csrfile_io_pageEn),
    .io_basePpn(csrfile_io_basePpn),
    .io_sum(csrfile_io_sum)
  );
  ExclusiveMonitor excMon ( // @[Core.scala 46:23]
    .clock(excMon_clock),
    .reset(excMon_reset),
    .io_flush(excMon_io_flush),
    .io_check_addr(excMon_io_check_addr),
    .io_check_valid(excMon_io_check_valid),
    .io_update_addr(excMon_io_update_addr),
    .io_update_set(excMon_io_update_set),
    .io_update_clear(excMon_io_update_clear)
  );
  HazardResolver resolve ( // @[Core.scala 49:23]
    .io_regRead1_en(resolve_io_regRead1_en),
    .io_regRead1_addr(resolve_io_regRead1_addr),
    .io_regRead1_data(resolve_io_regRead1_data),
    .io_regRead2_en(resolve_io_regRead2_en),
    .io_regRead2_addr(resolve_io_regRead2_addr),
    .io_regRead2_data(resolve_io_regRead2_data),
    .io_csrRead_op(resolve_io_csrRead_op),
    .io_csrRead_valid(resolve_io_csrRead_valid),
    .io_csrRead_addr(resolve_io_csrRead_addr),
    .io_csrRead_data(resolve_io_csrRead_data),
    .io_check_addr(resolve_io_check_addr),
    .io_check_valid(resolve_io_check_valid),
    .io_aluReg_en(resolve_io_aluReg_en),
    .io_aluReg_addr(resolve_io_aluReg_addr),
    .io_aluReg_data(resolve_io_aluReg_data),
    .io_aluReg_load(resolve_io_aluReg_load),
    .io_memReg_en(resolve_io_memReg_en),
    .io_memReg_addr(resolve_io_memReg_addr),
    .io_memReg_data(resolve_io_memReg_data),
    .io_memReg_load(resolve_io_memReg_load),
    .io_memCsr_op(resolve_io_memCsr_op),
    .io_memCsr_addr(resolve_io_memCsr_addr),
    .io_wbReg_en(resolve_io_wbReg_en),
    .io_wbReg_addr(resolve_io_wbReg_addr),
    .io_wbReg_data(resolve_io_wbReg_data),
    .io_wbCsr_op(resolve_io_wbCsr_op),
    .io_wbCsr_addr(resolve_io_wbCsr_addr),
    .io_wbExcMon_addr(resolve_io_wbExcMon_addr),
    .io_wbExcMon_set(resolve_io_wbExcMon_set),
    .io_wbExcMon_clear(resolve_io_wbExcMon_clear),
    .io_rf1_en(resolve_io_rf1_en),
    .io_rf1_addr(resolve_io_rf1_addr),
    .io_rf1_data(resolve_io_rf1_data),
    .io_rf2_en(resolve_io_rf2_en),
    .io_rf2_addr(resolve_io_rf2_addr),
    .io_rf2_data(resolve_io_rf2_data),
    .io_csr_op(resolve_io_csr_op),
    .io_csr_valid(resolve_io_csr_valid),
    .io_csr_addr(resolve_io_csr_addr),
    .io_csr_data(resolve_io_csr_data),
    .io_excMon_addr(resolve_io_excMon_addr),
    .io_excMon_valid(resolve_io_excMon_valid),
    .io_loadFlag(resolve_io_loadFlag),
    .io_csrFlag(resolve_io_csrFlag)
  );
  PipelineController control ( // @[Core.scala 50:23]
    .io_fetch(control_io_fetch),
    .io_alu(control_io_alu),
    .io_mem(control_io_mem),
    .io_decFlush(control_io_decFlush),
    .io_decTarget(control_io_decTarget),
    .io_memFlush(control_io_memFlush),
    .io_memTarget(control_io_memTarget),
    .io_load(control_io_load),
    .io_csr(control_io_csr),
    .io_except_hasTrap(control_io_except_hasTrap),
    .io_except_isSret(control_io_except_isSret),
    .io_except_isMret(control_io_except_isMret),
    .io_csrSepc(control_io_csrSepc),
    .io_csrMepc(control_io_csrMepc),
    .io_csrTvec(control_io_csrTvec),
    .io_stallIf(control_io_stallIf),
    .io_stallId(control_io_stallId),
    .io_stallEx(control_io_stallEx),
    .io_stallMm(control_io_stallMm),
    .io_stallWb(control_io_stallWb),
    .io_flush(control_io_flush),
    .io_flushIf(control_io_flushIf),
    .io_flushPc(control_io_flushPc)
  );
  assign io_tlb_en = csrfile_io_pageEn; // @[Core.scala 149:23]
  assign io_tlb_flushInst = mem_io_flushIt; // @[Core.scala 150:23]
  assign io_tlb_flushData = mem_io_flushDt; // @[Core.scala 151:23]
  assign io_tlb_basePpn = csrfile_io_basePpn; // @[Core.scala 152:23]
  assign io_tlb_sum = csrfile_io_sum; // @[Core.scala 153:23]
  assign io_tlb_smode = csrfile_io_mode[0]; // @[Core.scala 154:23]
  assign io_cache_flushInst = mem_io_flushIc; // @[Core.scala 155:23]
  assign io_cache_flushData = mem_io_flushDc; // @[Core.scala 156:23]
  assign io_rom_addr = fetch_io_rom_addr; // @[Core.scala 56:21]
  assign io_ram_en = mem_io_ram_en; // @[Core.scala 87:23]
  assign io_ram_wen = mem_io_ram_wen; // @[Core.scala 87:23]
  assign io_ram_addr = mem_io_ram_addr; // @[Core.scala 87:23]
  assign io_ram_wdata = mem_io_ram_wdata; // @[Core.scala 87:23]
  assign io_debug_regWen = wb_io_debug_regWen; // @[Core.scala 100:17]
  assign io_debug_regWaddr = wb_io_debug_regWaddr; // @[Core.scala 100:17]
  assign io_debug_regWdata = wb_io_debug_regWdata; // @[Core.scala 100:17]
  assign io_debug_pc = wb_io_debug_pc; // @[Core.scala 100:17]
  assign fetch_clock = clock;
  assign fetch_reset = reset;
  assign fetch_io_flush = control_io_flushIf; // @[Core.scala 53:21]
  assign fetch_io_stall = control_io_stallIf; // @[Core.scala 54:21]
  assign fetch_io_flushPc = control_io_flushPc; // @[Core.scala 55:21]
  assign fetch_io_rom_valid = io_rom_valid; // @[Core.scala 56:21]
  assign fetch_io_rom_fault = io_rom_fault; // @[Core.scala 56:21]
  assign fetch_io_branch_branch = decoder_io_branch_branch; // @[Core.scala 57:21]
  assign fetch_io_branch_jump = decoder_io_branch_jump; // @[Core.scala 57:21]
  assign fetch_io_branch_taken = decoder_io_branch_taken; // @[Core.scala 57:21]
  assign fetch_io_branch_index = decoder_io_branch_index; // @[Core.scala 57:21]
  assign fetch_io_branch_pc = decoder_io_branch_pc; // @[Core.scala 57:21]
  assign fetch_io_branch_target = decoder_io_branch_target; // @[Core.scala 57:21]
  assign ifid_clock = clock;
  assign ifid_reset = reset;
  assign ifid_io_flush = control_io_flushIf; // @[Core.scala 59:21]
  assign ifid_io_stallPrev = control_io_stallIf; // @[Core.scala 60:21]
  assign ifid_io_stallNext = control_io_stallId; // @[Core.scala 61:21]
  assign ifid_io_prev_valid = fetch_io_fetch_valid; // @[Core.scala 62:21]
  assign ifid_io_prev_pc = fetch_io_fetch_pc; // @[Core.scala 62:21]
  assign ifid_io_prev_taken = fetch_io_fetch_taken; // @[Core.scala 62:21]
  assign ifid_io_prev_target = fetch_io_fetch_target; // @[Core.scala 62:21]
  assign ifid_io_prev_predIndex = fetch_io_fetch_predIndex; // @[Core.scala 62:21]
  assign ifid_io_prev_pageFault = fetch_io_fetch_pageFault; // @[Core.scala 62:21]
  assign decoder_clock = clock;
  assign decoder_io_fetch_valid = ifid_io_next_valid; // @[Core.scala 65:23]
  assign decoder_io_fetch_pc = ifid_io_next_pc; // @[Core.scala 65:23]
  assign decoder_io_fetch_taken = ifid_io_next_taken; // @[Core.scala 65:23]
  assign decoder_io_fetch_target = ifid_io_next_target; // @[Core.scala 65:23]
  assign decoder_io_fetch_predIndex = ifid_io_next_predIndex; // @[Core.scala 65:23]
  assign decoder_io_fetch_pageFault = ifid_io_next_pageFault; // @[Core.scala 65:23]
  assign decoder_io_inst = io_rom_rdata; // @[Core.scala 66:23]
  assign decoder_io_stallId = control_io_stallId; // @[Core.scala 67:23]
  assign decoder_io_read1_data = resolve_io_regRead1_data; // @[Core.scala 68:23]
  assign decoder_io_read2_data = resolve_io_regRead2_data; // @[Core.scala 69:23]
  assign idex_clock = clock;
  assign idex_reset = reset;
  assign idex_io_flush = control_io_flush; // @[Core.scala 70:23]
  assign idex_io_stallPrev = control_io_stallId; // @[Core.scala 71:23]
  assign idex_io_stallNext = control_io_stallEx; // @[Core.scala 72:23]
  assign idex_io_prev_aluOp = decoder_io_decoder_aluOp; // @[Core.scala 73:23]
  assign idex_io_prev_opr1 = decoder_io_decoder_opr1; // @[Core.scala 73:23]
  assign idex_io_prev_opr2 = decoder_io_decoder_opr2; // @[Core.scala 73:23]
  assign idex_io_prev_mduOp = decoder_io_decoder_mduOp; // @[Core.scala 73:23]
  assign idex_io_prev_lsuOp = decoder_io_decoder_lsuOp; // @[Core.scala 73:23]
  assign idex_io_prev_lsuData = decoder_io_decoder_lsuData; // @[Core.scala 73:23]
  assign idex_io_prev_regWen = decoder_io_decoder_regWen; // @[Core.scala 73:23]
  assign idex_io_prev_regWaddr = decoder_io_decoder_regWaddr; // @[Core.scala 73:23]
  assign idex_io_prev_csrOp = decoder_io_decoder_csrOp; // @[Core.scala 73:23]
  assign idex_io_prev_csrAddr = decoder_io_decoder_csrAddr; // @[Core.scala 73:23]
  assign idex_io_prev_csrData = decoder_io_decoder_csrData; // @[Core.scala 73:23]
  assign idex_io_prev_excType = decoder_io_decoder_excType; // @[Core.scala 73:23]
  assign idex_io_prev_excValue = decoder_io_decoder_excValue; // @[Core.scala 73:23]
  assign idex_io_prev_valid = decoder_io_decoder_valid; // @[Core.scala 73:23]
  assign idex_io_prev_inst = decoder_io_decoder_inst; // @[Core.scala 73:23]
  assign idex_io_prev_currentPc = decoder_io_decoder_currentPc; // @[Core.scala 73:23]
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_decoder_aluOp = idex_io_next_aluOp; // @[Core.scala 76:23]
  assign alu_io_decoder_opr1 = idex_io_next_opr1; // @[Core.scala 76:23]
  assign alu_io_decoder_opr2 = idex_io_next_opr2; // @[Core.scala 76:23]
  assign alu_io_decoder_mduOp = idex_io_next_mduOp; // @[Core.scala 76:23]
  assign alu_io_decoder_lsuOp = idex_io_next_lsuOp; // @[Core.scala 76:23]
  assign alu_io_decoder_lsuData = idex_io_next_lsuData; // @[Core.scala 76:23]
  assign alu_io_decoder_regWen = idex_io_next_regWen; // @[Core.scala 76:23]
  assign alu_io_decoder_regWaddr = idex_io_next_regWaddr; // @[Core.scala 76:23]
  assign alu_io_decoder_csrOp = idex_io_next_csrOp; // @[Core.scala 76:23]
  assign alu_io_decoder_csrAddr = idex_io_next_csrAddr; // @[Core.scala 76:23]
  assign alu_io_decoder_csrData = idex_io_next_csrData; // @[Core.scala 76:23]
  assign alu_io_decoder_excType = idex_io_next_excType; // @[Core.scala 76:23]
  assign alu_io_decoder_excValue = idex_io_next_excValue; // @[Core.scala 76:23]
  assign alu_io_decoder_valid = idex_io_next_valid; // @[Core.scala 76:23]
  assign alu_io_decoder_inst = idex_io_next_inst; // @[Core.scala 76:23]
  assign alu_io_decoder_currentPc = idex_io_next_currentPc; // @[Core.scala 76:23]
  assign alu_io_flush = control_io_flush; // @[Core.scala 77:23]
  assign alu_io_csrRead_valid = resolve_io_csrRead_valid; // @[Core.scala 78:23]
  assign alu_io_csrRead_data = resolve_io_csrRead_data; // @[Core.scala 78:23]
  assign exmem_clock = clock;
  assign exmem_reset = reset;
  assign exmem_io_flush = control_io_flush; // @[Core.scala 79:23]
  assign exmem_io_stallPrev = control_io_stallEx; // @[Core.scala 80:23]
  assign exmem_io_stallNext = control_io_stallMm; // @[Core.scala 81:23]
  assign exmem_io_prev_lsuOp = alu_io_alu_lsuOp; // @[Core.scala 82:23]
  assign exmem_io_prev_lsuData = alu_io_alu_lsuData; // @[Core.scala 82:23]
  assign exmem_io_prev_reg_en = alu_io_alu_reg_en; // @[Core.scala 82:23]
  assign exmem_io_prev_reg_addr = alu_io_alu_reg_addr; // @[Core.scala 82:23]
  assign exmem_io_prev_reg_data = alu_io_alu_reg_data; // @[Core.scala 82:23]
  assign exmem_io_prev_csr_op = alu_io_alu_csr_op; // @[Core.scala 82:23]
  assign exmem_io_prev_csr_addr = alu_io_alu_csr_addr; // @[Core.scala 82:23]
  assign exmem_io_prev_csr_data = alu_io_alu_csr_data; // @[Core.scala 82:23]
  assign exmem_io_prev_csr_retired = alu_io_alu_csr_retired; // @[Core.scala 82:23]
  assign exmem_io_prev_excType = alu_io_alu_excType; // @[Core.scala 82:23]
  assign exmem_io_prev_excValue = alu_io_alu_excValue; // @[Core.scala 82:23]
  assign exmem_io_prev_valid = alu_io_alu_valid; // @[Core.scala 82:23]
  assign exmem_io_prev_inst = alu_io_alu_inst; // @[Core.scala 82:23]
  assign exmem_io_prev_currentPc = alu_io_alu_currentPc; // @[Core.scala 82:23]
  assign mem_clock = clock;
  assign mem_reset = reset;
  assign mem_io_alu_lsuOp = exmem_io_next_lsuOp; // @[Core.scala 85:23]
  assign mem_io_alu_lsuData = exmem_io_next_lsuData; // @[Core.scala 85:23]
  assign mem_io_alu_reg_en = exmem_io_next_reg_en; // @[Core.scala 85:23]
  assign mem_io_alu_reg_addr = exmem_io_next_reg_addr; // @[Core.scala 85:23]
  assign mem_io_alu_reg_data = exmem_io_next_reg_data; // @[Core.scala 85:23]
  assign mem_io_alu_csr_op = exmem_io_next_csr_op; // @[Core.scala 85:23]
  assign mem_io_alu_csr_addr = exmem_io_next_csr_addr; // @[Core.scala 85:23]
  assign mem_io_alu_csr_data = exmem_io_next_csr_data; // @[Core.scala 85:23]
  assign mem_io_alu_csr_retired = exmem_io_next_csr_retired; // @[Core.scala 85:23]
  assign mem_io_alu_excType = exmem_io_next_excType; // @[Core.scala 85:23]
  assign mem_io_alu_excValue = exmem_io_next_excValue; // @[Core.scala 85:23]
  assign mem_io_alu_valid = exmem_io_next_valid; // @[Core.scala 85:23]
  assign mem_io_alu_inst = exmem_io_next_inst; // @[Core.scala 85:23]
  assign mem_io_alu_currentPc = exmem_io_next_currentPc; // @[Core.scala 85:23]
  assign mem_io_flush = control_io_flush; // @[Core.scala 86:23]
  assign mem_io_ram_valid = io_ram_valid; // @[Core.scala 87:23]
  assign mem_io_ram_fault = io_ram_fault; // @[Core.scala 87:23]
  assign mem_io_ram_rdata = io_ram_rdata; // @[Core.scala 87:23]
  assign mem_io_csrHasInt = csrfile_io_hasInt; // @[Core.scala 88:23]
  assign mem_io_csrBusy = csrfile_io_busy; // @[Core.scala 89:23]
  assign mem_io_csrMode = csrfile_io_mode; // @[Core.scala 90:23]
  assign mem_io_excMon_valid = resolve_io_check_valid; // @[Core.scala 91:23]
  assign memwb_clock = clock;
  assign memwb_reset = reset;
  assign memwb_io_flush = control_io_flush; // @[Core.scala 92:23]
  assign memwb_io_stallPrev = control_io_stallMm; // @[Core.scala 93:23]
  assign memwb_io_stallNext = control_io_stallWb; // @[Core.scala 94:23]
  assign memwb_io_prev_reg_en = mem_io_mem_reg_en; // @[Core.scala 95:23]
  assign memwb_io_prev_reg_addr = mem_io_mem_reg_addr; // @[Core.scala 95:23]
  assign memwb_io_prev_reg_data = mem_io_mem_reg_data; // @[Core.scala 95:23]
  assign memwb_io_prev_reg_load = mem_io_mem_reg_load; // @[Core.scala 95:23]
  assign memwb_io_prev_memSigned = mem_io_mem_memSigned; // @[Core.scala 95:23]
  assign memwb_io_prev_memSel = mem_io_mem_memSel; // @[Core.scala 95:23]
  assign memwb_io_prev_memWidth = mem_io_mem_memWidth; // @[Core.scala 95:23]
  assign memwb_io_prev_csr_op = mem_io_mem_csr_op; // @[Core.scala 95:23]
  assign memwb_io_prev_csr_addr = mem_io_mem_csr_addr; // @[Core.scala 95:23]
  assign memwb_io_prev_csr_data = mem_io_mem_csr_data; // @[Core.scala 95:23]
  assign memwb_io_prev_csr_retired = mem_io_mem_csr_retired; // @[Core.scala 95:23]
  assign memwb_io_prev_excMon_addr = mem_io_mem_excMon_addr; // @[Core.scala 95:23]
  assign memwb_io_prev_excMon_set = mem_io_mem_excMon_set; // @[Core.scala 95:23]
  assign memwb_io_prev_excMon_clear = mem_io_mem_excMon_clear; // @[Core.scala 95:23]
  assign memwb_io_prev_currentPc = mem_io_mem_currentPc; // @[Core.scala 95:23]
  assign wb_io_mem_reg_en = memwb_io_next_reg_en; // @[Core.scala 98:17]
  assign wb_io_mem_reg_addr = memwb_io_next_reg_addr; // @[Core.scala 98:17]
  assign wb_io_mem_reg_data = memwb_io_next_reg_data; // @[Core.scala 98:17]
  assign wb_io_mem_reg_load = memwb_io_next_reg_load; // @[Core.scala 98:17]
  assign wb_io_mem_memSigned = memwb_io_next_memSigned; // @[Core.scala 98:17]
  assign wb_io_mem_memSel = memwb_io_next_memSel; // @[Core.scala 98:17]
  assign wb_io_mem_memWidth = memwb_io_next_memWidth; // @[Core.scala 98:17]
  assign wb_io_mem_csr_op = memwb_io_next_csr_op; // @[Core.scala 98:17]
  assign wb_io_mem_csr_addr = memwb_io_next_csr_addr; // @[Core.scala 98:17]
  assign wb_io_mem_csr_data = memwb_io_next_csr_data; // @[Core.scala 98:17]
  assign wb_io_mem_csr_retired = memwb_io_next_csr_retired; // @[Core.scala 98:17]
  assign wb_io_mem_excMon_addr = memwb_io_next_excMon_addr; // @[Core.scala 98:17]
  assign wb_io_mem_excMon_set = memwb_io_next_excMon_set; // @[Core.scala 98:17]
  assign wb_io_mem_excMon_clear = memwb_io_next_excMon_clear; // @[Core.scala 98:17]
  assign wb_io_mem_currentPc = memwb_io_next_currentPc; // @[Core.scala 98:17]
  assign wb_io_ramData = io_ram_rdata; // @[Core.scala 99:17]
  assign regfile_clock = clock;
  assign regfile_reset = reset;
  assign regfile_io_read1_en = resolve_io_rf1_en; // @[Core.scala 103:25]
  assign regfile_io_read1_addr = resolve_io_rf1_addr; // @[Core.scala 103:25]
  assign regfile_io_read2_en = resolve_io_rf2_en; // @[Core.scala 104:25]
  assign regfile_io_read2_addr = resolve_io_rf2_addr; // @[Core.scala 104:25]
  assign regfile_io_write_en = wb_io_reg_en; // @[Core.scala 105:25]
  assign regfile_io_write_addr = wb_io_reg_addr; // @[Core.scala 106:25]
  assign regfile_io_write_data = wb_io_reg_data; // @[Core.scala 107:25]
  assign csrfile_clock = clock;
  assign csrfile_reset = reset;
  assign csrfile_io_read_op = resolve_io_csr_op; // @[Core.scala 110:29]
  assign csrfile_io_read_addr = resolve_io_csr_addr; // @[Core.scala 110:29]
  assign csrfile_io_write_op = wb_io_csr_op; // @[Core.scala 111:29]
  assign csrfile_io_write_addr = wb_io_csr_addr; // @[Core.scala 112:29]
  assign csrfile_io_write_data = wb_io_csr_data; // @[Core.scala 113:29]
  assign csrfile_io_write_retired = wb_io_csr_retired; // @[Core.scala 114:29]
  assign csrfile_io_irq_timer = io_irq_timer; // @[Core.scala 115:29]
  assign csrfile_io_irq_soft = io_irq_soft; // @[Core.scala 115:29]
  assign csrfile_io_irq_extern = io_irq_extern; // @[Core.scala 115:29]
  assign csrfile_io_except_hasTrap = mem_io_except_hasTrap; // @[Core.scala 116:29]
  assign csrfile_io_except_isSret = mem_io_except_isSret; // @[Core.scala 116:29]
  assign csrfile_io_except_isMret = mem_io_except_isMret; // @[Core.scala 116:29]
  assign csrfile_io_except_excCause = mem_io_except_excCause; // @[Core.scala 116:29]
  assign csrfile_io_except_excPc = mem_io_except_excPc; // @[Core.scala 116:29]
  assign csrfile_io_except_excValue = mem_io_except_excValue; // @[Core.scala 116:29]
  assign excMon_clock = clock;
  assign excMon_reset = reset;
  assign excMon_io_flush = control_io_flush; // @[Core.scala 119:27]
  assign excMon_io_check_addr = resolve_io_excMon_addr; // @[Core.scala 120:27]
  assign excMon_io_update_addr = wb_io_excMon_addr; // @[Core.scala 121:27]
  assign excMon_io_update_set = wb_io_excMon_set; // @[Core.scala 122:27]
  assign excMon_io_update_clear = wb_io_excMon_clear; // @[Core.scala 123:27]
  assign resolve_io_regRead1_en = decoder_io_read1_en; // @[Core.scala 68:23]
  assign resolve_io_regRead1_addr = decoder_io_read1_addr; // @[Core.scala 68:23]
  assign resolve_io_regRead2_en = decoder_io_read2_en; // @[Core.scala 69:23]
  assign resolve_io_regRead2_addr = decoder_io_read2_addr; // @[Core.scala 69:23]
  assign resolve_io_csrRead_op = alu_io_csrRead_op; // @[Core.scala 78:23]
  assign resolve_io_csrRead_addr = alu_io_csrRead_addr; // @[Core.scala 78:23]
  assign resolve_io_check_addr = mem_io_excMon_addr; // @[Core.scala 91:23]
  assign resolve_io_aluReg_en = alu_io_alu_reg_en; // @[Core.scala 126:23]
  assign resolve_io_aluReg_addr = alu_io_alu_reg_addr; // @[Core.scala 126:23]
  assign resolve_io_aluReg_data = alu_io_alu_reg_data; // @[Core.scala 126:23]
  assign resolve_io_aluReg_load = alu_io_alu_reg_load; // @[Core.scala 126:23]
  assign resolve_io_memReg_en = mem_io_mem_reg_en; // @[Core.scala 127:23]
  assign resolve_io_memReg_addr = mem_io_mem_reg_addr; // @[Core.scala 127:23]
  assign resolve_io_memReg_data = mem_io_mem_reg_data; // @[Core.scala 127:23]
  assign resolve_io_memReg_load = mem_io_mem_reg_load; // @[Core.scala 127:23]
  assign resolve_io_memCsr_op = mem_io_mem_csr_op; // @[Core.scala 128:23]
  assign resolve_io_memCsr_addr = mem_io_mem_csr_addr; // @[Core.scala 128:23]
  assign resolve_io_wbReg_en = wb_io_reg_en; // @[Core.scala 129:23]
  assign resolve_io_wbReg_addr = wb_io_reg_addr; // @[Core.scala 129:23]
  assign resolve_io_wbReg_data = wb_io_reg_data; // @[Core.scala 129:23]
  assign resolve_io_wbCsr_op = wb_io_csr_op; // @[Core.scala 130:23]
  assign resolve_io_wbCsr_addr = wb_io_csr_addr; // @[Core.scala 130:23]
  assign resolve_io_wbExcMon_addr = wb_io_excMon_addr; // @[Core.scala 131:23]
  assign resolve_io_wbExcMon_set = wb_io_excMon_set; // @[Core.scala 131:23]
  assign resolve_io_wbExcMon_clear = wb_io_excMon_clear; // @[Core.scala 131:23]
  assign resolve_io_rf1_data = regfile_io_read1_data; // @[Core.scala 103:25]
  assign resolve_io_rf2_data = regfile_io_read2_data; // @[Core.scala 104:25]
  assign resolve_io_csr_valid = csrfile_io_read_valid; // @[Core.scala 110:29]
  assign resolve_io_csr_data = csrfile_io_read_data; // @[Core.scala 110:29]
  assign resolve_io_excMon_valid = excMon_io_check_valid; // @[Core.scala 120:27]
  assign control_io_fetch = fetch_io_stallReq; // @[Core.scala 134:25]
  assign control_io_alu = alu_io_stallReq; // @[Core.scala 135:25]
  assign control_io_mem = mem_io_stallReq; // @[Core.scala 136:25]
  assign control_io_decFlush = decoder_io_flushIf; // @[Core.scala 137:25]
  assign control_io_decTarget = decoder_io_flushPc; // @[Core.scala 138:25]
  assign control_io_memFlush = mem_io_flushReq; // @[Core.scala 139:25]
  assign control_io_memTarget = mem_io_flushPc; // @[Core.scala 140:25]
  assign control_io_load = resolve_io_loadFlag; // @[Core.scala 141:25]
  assign control_io_csr = resolve_io_csrFlag; // @[Core.scala 142:25]
  assign control_io_except_hasTrap = mem_io_except_hasTrap; // @[Core.scala 143:25]
  assign control_io_except_isSret = mem_io_except_isSret; // @[Core.scala 143:25]
  assign control_io_except_isMret = mem_io_except_isMret; // @[Core.scala 143:25]
  assign control_io_csrSepc = csrfile_io_sepc; // @[Core.scala 144:25]
  assign control_io_csrMepc = csrfile_io_mepc; // @[Core.scala 145:25]
  assign control_io_csrTvec = csrfile_io_trapVec; // @[Core.scala 146:25]
endmodule
module TLB(
  input         clock,
  input         reset,
  input         io_flush,
  input         io_wen,
  input  [31:0] io_vaddr,
  input  [21:0] io_went_ppn,
  input         io_went_d,
  input         io_went_a,
  input         io_went_u,
  input         io_went_x,
  input         io_went_w,
  input         io_went_r,
  output        io_valid,
  output [21:0] io_rent_ppn,
  output        io_rent_d,
  output        io_rent_a,
  output        io_rent_u,
  output        io_rent_x,
  output        io_rent_w,
  output        io_rent_r
);
  reg [19:0] data_vpn [0:15]; // @[TLB.scala 37:18]
  reg [31:0] _RAND_0;
  wire [19:0] data_vpn__T_6_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_6_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_9_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_9_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_10_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_10_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_13_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_13_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_14_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_14_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_17_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_17_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_18_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_18_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_21_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_21_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_22_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_22_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_25_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_25_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_26_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_26_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_29_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_29_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_30_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_30_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_33_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_33_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_34_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_34_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_37_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_37_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_38_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_38_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_41_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_41_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_42_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_42_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_45_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_45_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_46_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_46_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_49_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_49_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_50_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_50_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_53_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_53_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_54_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_54_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_57_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_57_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_58_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_58_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_61_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_61_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_62_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_62_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_65_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_65_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_66_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_66_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_69_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_69_addr; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_1_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_1_addr; // @[TLB.scala 37:18]
  wire  data_vpn__T_1_mask; // @[TLB.scala 37:18]
  wire  data_vpn__T_1_en; // @[TLB.scala 37:18]
  wire [19:0] data_vpn__T_2_data; // @[TLB.scala 37:18]
  wire [3:0] data_vpn__T_2_addr; // @[TLB.scala 37:18]
  wire  data_vpn__T_2_mask; // @[TLB.scala 37:18]
  wire  data_vpn__T_2_en; // @[TLB.scala 37:18]
  reg [21:0] data_entry_ppn [0:15]; // @[TLB.scala 37:18]
  reg [31:0] _RAND_1;
  wire [21:0] data_entry_ppn__T_6_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_6_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_9_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_9_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_10_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_10_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_13_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_13_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_14_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_14_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_17_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_17_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_18_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_18_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_21_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_21_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_22_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_22_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_25_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_25_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_26_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_26_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_29_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_29_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_30_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_30_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_33_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_33_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_34_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_34_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_37_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_37_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_38_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_38_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_41_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_41_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_42_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_42_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_45_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_45_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_46_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_46_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_49_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_49_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_50_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_50_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_53_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_53_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_54_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_54_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_57_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_57_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_58_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_58_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_61_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_61_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_62_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_62_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_65_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_65_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_66_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_66_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_69_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_69_addr; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_1_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_1_addr; // @[TLB.scala 37:18]
  wire  data_entry_ppn__T_1_mask; // @[TLB.scala 37:18]
  wire  data_entry_ppn__T_1_en; // @[TLB.scala 37:18]
  wire [21:0] data_entry_ppn__T_2_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_ppn__T_2_addr; // @[TLB.scala 37:18]
  wire  data_entry_ppn__T_2_mask; // @[TLB.scala 37:18]
  wire  data_entry_ppn__T_2_en; // @[TLB.scala 37:18]
  reg  data_entry_d [0:15]; // @[TLB.scala 37:18]
  reg [31:0] _RAND_2;
  wire  data_entry_d__T_6_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_6_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_9_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_9_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_10_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_10_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_13_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_13_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_14_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_14_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_17_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_17_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_18_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_18_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_21_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_21_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_22_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_22_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_25_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_25_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_26_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_26_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_29_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_29_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_30_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_30_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_33_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_33_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_34_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_34_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_37_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_37_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_38_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_38_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_41_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_41_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_42_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_42_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_45_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_45_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_46_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_46_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_49_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_49_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_50_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_50_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_53_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_53_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_54_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_54_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_57_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_57_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_58_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_58_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_61_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_61_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_62_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_62_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_65_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_65_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_66_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_66_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_69_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_69_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_1_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_1_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_1_mask; // @[TLB.scala 37:18]
  wire  data_entry_d__T_1_en; // @[TLB.scala 37:18]
  wire  data_entry_d__T_2_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_d__T_2_addr; // @[TLB.scala 37:18]
  wire  data_entry_d__T_2_mask; // @[TLB.scala 37:18]
  wire  data_entry_d__T_2_en; // @[TLB.scala 37:18]
  reg  data_entry_a [0:15]; // @[TLB.scala 37:18]
  reg [31:0] _RAND_3;
  wire  data_entry_a__T_6_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_6_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_9_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_9_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_10_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_10_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_13_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_13_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_14_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_14_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_17_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_17_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_18_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_18_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_21_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_21_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_22_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_22_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_25_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_25_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_26_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_26_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_29_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_29_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_30_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_30_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_33_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_33_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_34_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_34_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_37_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_37_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_38_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_38_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_41_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_41_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_42_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_42_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_45_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_45_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_46_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_46_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_49_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_49_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_50_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_50_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_53_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_53_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_54_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_54_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_57_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_57_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_58_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_58_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_61_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_61_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_62_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_62_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_65_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_65_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_66_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_66_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_69_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_69_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_1_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_1_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_1_mask; // @[TLB.scala 37:18]
  wire  data_entry_a__T_1_en; // @[TLB.scala 37:18]
  wire  data_entry_a__T_2_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_a__T_2_addr; // @[TLB.scala 37:18]
  wire  data_entry_a__T_2_mask; // @[TLB.scala 37:18]
  wire  data_entry_a__T_2_en; // @[TLB.scala 37:18]
  reg  data_entry_u [0:15]; // @[TLB.scala 37:18]
  reg [31:0] _RAND_4;
  wire  data_entry_u__T_6_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_6_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_9_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_9_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_10_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_10_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_13_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_13_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_14_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_14_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_17_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_17_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_18_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_18_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_21_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_21_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_22_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_22_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_25_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_25_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_26_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_26_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_29_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_29_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_30_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_30_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_33_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_33_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_34_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_34_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_37_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_37_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_38_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_38_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_41_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_41_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_42_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_42_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_45_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_45_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_46_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_46_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_49_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_49_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_50_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_50_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_53_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_53_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_54_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_54_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_57_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_57_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_58_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_58_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_61_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_61_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_62_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_62_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_65_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_65_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_66_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_66_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_69_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_69_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_1_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_1_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_1_mask; // @[TLB.scala 37:18]
  wire  data_entry_u__T_1_en; // @[TLB.scala 37:18]
  wire  data_entry_u__T_2_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_u__T_2_addr; // @[TLB.scala 37:18]
  wire  data_entry_u__T_2_mask; // @[TLB.scala 37:18]
  wire  data_entry_u__T_2_en; // @[TLB.scala 37:18]
  reg  data_entry_x [0:15]; // @[TLB.scala 37:18]
  reg [31:0] _RAND_5;
  wire  data_entry_x__T_6_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_6_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_9_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_9_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_10_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_10_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_13_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_13_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_14_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_14_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_17_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_17_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_18_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_18_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_21_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_21_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_22_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_22_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_25_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_25_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_26_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_26_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_29_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_29_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_30_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_30_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_33_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_33_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_34_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_34_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_37_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_37_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_38_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_38_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_41_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_41_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_42_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_42_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_45_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_45_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_46_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_46_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_49_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_49_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_50_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_50_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_53_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_53_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_54_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_54_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_57_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_57_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_58_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_58_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_61_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_61_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_62_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_62_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_65_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_65_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_66_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_66_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_69_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_69_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_1_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_1_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_1_mask; // @[TLB.scala 37:18]
  wire  data_entry_x__T_1_en; // @[TLB.scala 37:18]
  wire  data_entry_x__T_2_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_x__T_2_addr; // @[TLB.scala 37:18]
  wire  data_entry_x__T_2_mask; // @[TLB.scala 37:18]
  wire  data_entry_x__T_2_en; // @[TLB.scala 37:18]
  reg  data_entry_w [0:15]; // @[TLB.scala 37:18]
  reg [31:0] _RAND_6;
  wire  data_entry_w__T_6_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_6_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_9_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_9_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_10_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_10_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_13_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_13_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_14_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_14_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_17_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_17_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_18_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_18_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_21_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_21_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_22_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_22_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_25_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_25_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_26_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_26_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_29_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_29_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_30_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_30_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_33_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_33_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_34_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_34_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_37_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_37_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_38_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_38_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_41_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_41_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_42_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_42_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_45_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_45_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_46_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_46_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_49_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_49_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_50_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_50_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_53_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_53_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_54_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_54_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_57_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_57_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_58_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_58_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_61_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_61_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_62_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_62_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_65_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_65_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_66_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_66_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_69_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_69_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_1_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_1_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_1_mask; // @[TLB.scala 37:18]
  wire  data_entry_w__T_1_en; // @[TLB.scala 37:18]
  wire  data_entry_w__T_2_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_w__T_2_addr; // @[TLB.scala 37:18]
  wire  data_entry_w__T_2_mask; // @[TLB.scala 37:18]
  wire  data_entry_w__T_2_en; // @[TLB.scala 37:18]
  reg  data_entry_r [0:15]; // @[TLB.scala 37:18]
  reg [31:0] _RAND_7;
  wire  data_entry_r__T_6_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_6_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_9_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_9_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_10_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_10_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_13_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_13_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_14_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_14_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_17_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_17_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_18_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_18_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_21_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_21_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_22_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_22_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_25_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_25_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_26_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_26_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_29_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_29_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_30_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_30_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_33_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_33_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_34_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_34_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_37_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_37_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_38_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_38_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_41_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_41_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_42_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_42_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_45_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_45_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_46_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_46_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_49_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_49_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_50_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_50_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_53_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_53_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_54_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_54_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_57_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_57_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_58_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_58_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_61_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_61_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_62_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_62_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_65_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_65_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_66_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_66_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_69_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_69_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_1_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_1_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_1_mask; // @[TLB.scala 37:18]
  wire  data_entry_r__T_1_en; // @[TLB.scala 37:18]
  wire  data_entry_r__T_2_data; // @[TLB.scala 37:18]
  wire [3:0] data_entry_r__T_2_addr; // @[TLB.scala 37:18]
  wire  data_entry_r__T_2_mask; // @[TLB.scala 37:18]
  wire  data_entry_r__T_2_en; // @[TLB.scala 37:18]
  reg  valid_0; // @[TLB.scala 36:22]
  reg [31:0] _RAND_8;
  reg  valid_1; // @[TLB.scala 36:22]
  reg [31:0] _RAND_9;
  reg  valid_2; // @[TLB.scala 36:22]
  reg [31:0] _RAND_10;
  reg  valid_3; // @[TLB.scala 36:22]
  reg [31:0] _RAND_11;
  reg  valid_4; // @[TLB.scala 36:22]
  reg [31:0] _RAND_12;
  reg  valid_5; // @[TLB.scala 36:22]
  reg [31:0] _RAND_13;
  reg  valid_6; // @[TLB.scala 36:22]
  reg [31:0] _RAND_14;
  reg  valid_7; // @[TLB.scala 36:22]
  reg [31:0] _RAND_15;
  reg  valid_8; // @[TLB.scala 36:22]
  reg [31:0] _RAND_16;
  reg  valid_9; // @[TLB.scala 36:22]
  reg [31:0] _RAND_17;
  reg  valid_10; // @[TLB.scala 36:22]
  reg [31:0] _RAND_18;
  reg  valid_11; // @[TLB.scala 36:22]
  reg [31:0] _RAND_19;
  reg  valid_12; // @[TLB.scala 36:22]
  reg [31:0] _RAND_20;
  reg  valid_13; // @[TLB.scala 36:22]
  reg [31:0] _RAND_21;
  reg  valid_14; // @[TLB.scala 36:22]
  reg [31:0] _RAND_22;
  reg  valid_15; // @[TLB.scala 36:22]
  reg [31:0] _RAND_23;
  reg [3:0] pointer; // @[TLB.scala 43:24]
  reg [31:0] _RAND_24;
  wire [19:0] vpn = io_vaddr[31:12]; // @[TLB.scala 44:25]
  wire  _GEN_251 = 4'h0 == pointer; // @[TLB.scala 52:25]
  wire  _GEN_0 = _GEN_251 | valid_0; // @[TLB.scala 52:25]
  wire  _GEN_252 = 4'h1 == pointer; // @[TLB.scala 52:25]
  wire  _GEN_1 = _GEN_252 | valid_1; // @[TLB.scala 52:25]
  wire  _GEN_253 = 4'h2 == pointer; // @[TLB.scala 52:25]
  wire  _GEN_2 = _GEN_253 | valid_2; // @[TLB.scala 52:25]
  wire  _GEN_254 = 4'h3 == pointer; // @[TLB.scala 52:25]
  wire  _GEN_3 = _GEN_254 | valid_3; // @[TLB.scala 52:25]
  wire  _GEN_255 = 4'h4 == pointer; // @[TLB.scala 52:25]
  wire  _GEN_4 = _GEN_255 | valid_4; // @[TLB.scala 52:25]
  wire  _GEN_256 = 4'h5 == pointer; // @[TLB.scala 52:25]
  wire  _GEN_5 = _GEN_256 | valid_5; // @[TLB.scala 52:25]
  wire  _GEN_257 = 4'h6 == pointer; // @[TLB.scala 52:25]
  wire  _GEN_6 = _GEN_257 | valid_6; // @[TLB.scala 52:25]
  wire  _GEN_258 = 4'h7 == pointer; // @[TLB.scala 52:25]
  wire  _GEN_7 = _GEN_258 | valid_7; // @[TLB.scala 52:25]
  wire  _GEN_259 = 4'h8 == pointer; // @[TLB.scala 52:25]
  wire  _GEN_8 = _GEN_259 | valid_8; // @[TLB.scala 52:25]
  wire  _GEN_260 = 4'h9 == pointer; // @[TLB.scala 52:25]
  wire  _GEN_9 = _GEN_260 | valid_9; // @[TLB.scala 52:25]
  wire  _GEN_261 = 4'ha == pointer; // @[TLB.scala 52:25]
  wire  _GEN_10 = _GEN_261 | valid_10; // @[TLB.scala 52:25]
  wire  _GEN_262 = 4'hb == pointer; // @[TLB.scala 52:25]
  wire  _GEN_11 = _GEN_262 | valid_11; // @[TLB.scala 52:25]
  wire  _GEN_263 = 4'hc == pointer; // @[TLB.scala 52:25]
  wire  _GEN_12 = _GEN_263 | valid_12; // @[TLB.scala 52:25]
  wire  _GEN_264 = 4'hd == pointer; // @[TLB.scala 52:25]
  wire  _GEN_13 = _GEN_264 | valid_13; // @[TLB.scala 52:25]
  wire  _GEN_265 = 4'he == pointer; // @[TLB.scala 52:25]
  wire  _GEN_14 = _GEN_265 | valid_14; // @[TLB.scala 52:25]
  wire  _GEN_266 = 4'hf == pointer; // @[TLB.scala 52:25]
  wire  _GEN_15 = _GEN_266 | valid_15; // @[TLB.scala 52:25]
  wire [3:0] _T_4 = pointer + 4'h1; // @[TLB.scala 56:24]
  wire  _T_7 = data_vpn__T_6_data == vpn; // @[TLB.scala 63:35]
  wire  _T_8 = valid_0 & _T_7; // @[TLB.scala 63:20]
  wire  _GEN_79 = _T_8 & data_entry_r__T_9_data; // @[TLB.scala 63:44]
  wire  _GEN_80 = _T_8 & data_entry_w__T_9_data; // @[TLB.scala 63:44]
  wire  _GEN_81 = _T_8 & data_entry_x__T_9_data; // @[TLB.scala 63:44]
  wire  _GEN_82 = _T_8 & data_entry_u__T_9_data; // @[TLB.scala 63:44]
  wire  _GEN_83 = _T_8 & data_entry_a__T_9_data; // @[TLB.scala 63:44]
  wire  _GEN_84 = _T_8 & data_entry_d__T_9_data; // @[TLB.scala 63:44]
  wire [21:0] _GEN_85 = _T_8 ? data_entry_ppn__T_9_data : 22'h0; // @[TLB.scala 63:44]
  wire  _T_11 = data_vpn__T_10_data == vpn; // @[TLB.scala 63:35]
  wire  _T_12 = valid_1 & _T_11; // @[TLB.scala 63:20]
  wire  _GEN_86 = _T_12 | _T_8; // @[TLB.scala 63:44]
  wire  _GEN_90 = _T_12 ? data_entry_r__T_13_data : _GEN_79; // @[TLB.scala 63:44]
  wire  _GEN_91 = _T_12 ? data_entry_w__T_13_data : _GEN_80; // @[TLB.scala 63:44]
  wire  _GEN_92 = _T_12 ? data_entry_x__T_13_data : _GEN_81; // @[TLB.scala 63:44]
  wire  _GEN_93 = _T_12 ? data_entry_u__T_13_data : _GEN_82; // @[TLB.scala 63:44]
  wire  _GEN_94 = _T_12 ? data_entry_a__T_13_data : _GEN_83; // @[TLB.scala 63:44]
  wire  _GEN_95 = _T_12 ? data_entry_d__T_13_data : _GEN_84; // @[TLB.scala 63:44]
  wire [21:0] _GEN_96 = _T_12 ? data_entry_ppn__T_13_data : _GEN_85; // @[TLB.scala 63:44]
  wire  _T_15 = data_vpn__T_14_data == vpn; // @[TLB.scala 63:35]
  wire  _T_16 = valid_2 & _T_15; // @[TLB.scala 63:20]
  wire  _GEN_97 = _T_16 | _GEN_86; // @[TLB.scala 63:44]
  wire  _GEN_101 = _T_16 ? data_entry_r__T_17_data : _GEN_90; // @[TLB.scala 63:44]
  wire  _GEN_102 = _T_16 ? data_entry_w__T_17_data : _GEN_91; // @[TLB.scala 63:44]
  wire  _GEN_103 = _T_16 ? data_entry_x__T_17_data : _GEN_92; // @[TLB.scala 63:44]
  wire  _GEN_104 = _T_16 ? data_entry_u__T_17_data : _GEN_93; // @[TLB.scala 63:44]
  wire  _GEN_105 = _T_16 ? data_entry_a__T_17_data : _GEN_94; // @[TLB.scala 63:44]
  wire  _GEN_106 = _T_16 ? data_entry_d__T_17_data : _GEN_95; // @[TLB.scala 63:44]
  wire [21:0] _GEN_107 = _T_16 ? data_entry_ppn__T_17_data : _GEN_96; // @[TLB.scala 63:44]
  wire  _T_19 = data_vpn__T_18_data == vpn; // @[TLB.scala 63:35]
  wire  _T_20 = valid_3 & _T_19; // @[TLB.scala 63:20]
  wire  _GEN_108 = _T_20 | _GEN_97; // @[TLB.scala 63:44]
  wire  _GEN_112 = _T_20 ? data_entry_r__T_21_data : _GEN_101; // @[TLB.scala 63:44]
  wire  _GEN_113 = _T_20 ? data_entry_w__T_21_data : _GEN_102; // @[TLB.scala 63:44]
  wire  _GEN_114 = _T_20 ? data_entry_x__T_21_data : _GEN_103; // @[TLB.scala 63:44]
  wire  _GEN_115 = _T_20 ? data_entry_u__T_21_data : _GEN_104; // @[TLB.scala 63:44]
  wire  _GEN_116 = _T_20 ? data_entry_a__T_21_data : _GEN_105; // @[TLB.scala 63:44]
  wire  _GEN_117 = _T_20 ? data_entry_d__T_21_data : _GEN_106; // @[TLB.scala 63:44]
  wire [21:0] _GEN_118 = _T_20 ? data_entry_ppn__T_21_data : _GEN_107; // @[TLB.scala 63:44]
  wire  _T_23 = data_vpn__T_22_data == vpn; // @[TLB.scala 63:35]
  wire  _T_24 = valid_4 & _T_23; // @[TLB.scala 63:20]
  wire  _GEN_119 = _T_24 | _GEN_108; // @[TLB.scala 63:44]
  wire  _GEN_123 = _T_24 ? data_entry_r__T_25_data : _GEN_112; // @[TLB.scala 63:44]
  wire  _GEN_124 = _T_24 ? data_entry_w__T_25_data : _GEN_113; // @[TLB.scala 63:44]
  wire  _GEN_125 = _T_24 ? data_entry_x__T_25_data : _GEN_114; // @[TLB.scala 63:44]
  wire  _GEN_126 = _T_24 ? data_entry_u__T_25_data : _GEN_115; // @[TLB.scala 63:44]
  wire  _GEN_127 = _T_24 ? data_entry_a__T_25_data : _GEN_116; // @[TLB.scala 63:44]
  wire  _GEN_128 = _T_24 ? data_entry_d__T_25_data : _GEN_117; // @[TLB.scala 63:44]
  wire [21:0] _GEN_129 = _T_24 ? data_entry_ppn__T_25_data : _GEN_118; // @[TLB.scala 63:44]
  wire  _T_27 = data_vpn__T_26_data == vpn; // @[TLB.scala 63:35]
  wire  _T_28 = valid_5 & _T_27; // @[TLB.scala 63:20]
  wire  _GEN_130 = _T_28 | _GEN_119; // @[TLB.scala 63:44]
  wire  _GEN_134 = _T_28 ? data_entry_r__T_29_data : _GEN_123; // @[TLB.scala 63:44]
  wire  _GEN_135 = _T_28 ? data_entry_w__T_29_data : _GEN_124; // @[TLB.scala 63:44]
  wire  _GEN_136 = _T_28 ? data_entry_x__T_29_data : _GEN_125; // @[TLB.scala 63:44]
  wire  _GEN_137 = _T_28 ? data_entry_u__T_29_data : _GEN_126; // @[TLB.scala 63:44]
  wire  _GEN_138 = _T_28 ? data_entry_a__T_29_data : _GEN_127; // @[TLB.scala 63:44]
  wire  _GEN_139 = _T_28 ? data_entry_d__T_29_data : _GEN_128; // @[TLB.scala 63:44]
  wire [21:0] _GEN_140 = _T_28 ? data_entry_ppn__T_29_data : _GEN_129; // @[TLB.scala 63:44]
  wire  _T_31 = data_vpn__T_30_data == vpn; // @[TLB.scala 63:35]
  wire  _T_32 = valid_6 & _T_31; // @[TLB.scala 63:20]
  wire  _GEN_141 = _T_32 | _GEN_130; // @[TLB.scala 63:44]
  wire  _GEN_145 = _T_32 ? data_entry_r__T_33_data : _GEN_134; // @[TLB.scala 63:44]
  wire  _GEN_146 = _T_32 ? data_entry_w__T_33_data : _GEN_135; // @[TLB.scala 63:44]
  wire  _GEN_147 = _T_32 ? data_entry_x__T_33_data : _GEN_136; // @[TLB.scala 63:44]
  wire  _GEN_148 = _T_32 ? data_entry_u__T_33_data : _GEN_137; // @[TLB.scala 63:44]
  wire  _GEN_149 = _T_32 ? data_entry_a__T_33_data : _GEN_138; // @[TLB.scala 63:44]
  wire  _GEN_150 = _T_32 ? data_entry_d__T_33_data : _GEN_139; // @[TLB.scala 63:44]
  wire [21:0] _GEN_151 = _T_32 ? data_entry_ppn__T_33_data : _GEN_140; // @[TLB.scala 63:44]
  wire  _T_35 = data_vpn__T_34_data == vpn; // @[TLB.scala 63:35]
  wire  _T_36 = valid_7 & _T_35; // @[TLB.scala 63:20]
  wire  _GEN_152 = _T_36 | _GEN_141; // @[TLB.scala 63:44]
  wire  _GEN_156 = _T_36 ? data_entry_r__T_37_data : _GEN_145; // @[TLB.scala 63:44]
  wire  _GEN_157 = _T_36 ? data_entry_w__T_37_data : _GEN_146; // @[TLB.scala 63:44]
  wire  _GEN_158 = _T_36 ? data_entry_x__T_37_data : _GEN_147; // @[TLB.scala 63:44]
  wire  _GEN_159 = _T_36 ? data_entry_u__T_37_data : _GEN_148; // @[TLB.scala 63:44]
  wire  _GEN_160 = _T_36 ? data_entry_a__T_37_data : _GEN_149; // @[TLB.scala 63:44]
  wire  _GEN_161 = _T_36 ? data_entry_d__T_37_data : _GEN_150; // @[TLB.scala 63:44]
  wire [21:0] _GEN_162 = _T_36 ? data_entry_ppn__T_37_data : _GEN_151; // @[TLB.scala 63:44]
  wire  _T_39 = data_vpn__T_38_data == vpn; // @[TLB.scala 63:35]
  wire  _T_40 = valid_8 & _T_39; // @[TLB.scala 63:20]
  wire  _GEN_163 = _T_40 | _GEN_152; // @[TLB.scala 63:44]
  wire  _GEN_167 = _T_40 ? data_entry_r__T_41_data : _GEN_156; // @[TLB.scala 63:44]
  wire  _GEN_168 = _T_40 ? data_entry_w__T_41_data : _GEN_157; // @[TLB.scala 63:44]
  wire  _GEN_169 = _T_40 ? data_entry_x__T_41_data : _GEN_158; // @[TLB.scala 63:44]
  wire  _GEN_170 = _T_40 ? data_entry_u__T_41_data : _GEN_159; // @[TLB.scala 63:44]
  wire  _GEN_171 = _T_40 ? data_entry_a__T_41_data : _GEN_160; // @[TLB.scala 63:44]
  wire  _GEN_172 = _T_40 ? data_entry_d__T_41_data : _GEN_161; // @[TLB.scala 63:44]
  wire [21:0] _GEN_173 = _T_40 ? data_entry_ppn__T_41_data : _GEN_162; // @[TLB.scala 63:44]
  wire  _T_43 = data_vpn__T_42_data == vpn; // @[TLB.scala 63:35]
  wire  _T_44 = valid_9 & _T_43; // @[TLB.scala 63:20]
  wire  _GEN_174 = _T_44 | _GEN_163; // @[TLB.scala 63:44]
  wire  _GEN_178 = _T_44 ? data_entry_r__T_45_data : _GEN_167; // @[TLB.scala 63:44]
  wire  _GEN_179 = _T_44 ? data_entry_w__T_45_data : _GEN_168; // @[TLB.scala 63:44]
  wire  _GEN_180 = _T_44 ? data_entry_x__T_45_data : _GEN_169; // @[TLB.scala 63:44]
  wire  _GEN_181 = _T_44 ? data_entry_u__T_45_data : _GEN_170; // @[TLB.scala 63:44]
  wire  _GEN_182 = _T_44 ? data_entry_a__T_45_data : _GEN_171; // @[TLB.scala 63:44]
  wire  _GEN_183 = _T_44 ? data_entry_d__T_45_data : _GEN_172; // @[TLB.scala 63:44]
  wire [21:0] _GEN_184 = _T_44 ? data_entry_ppn__T_45_data : _GEN_173; // @[TLB.scala 63:44]
  wire  _T_47 = data_vpn__T_46_data == vpn; // @[TLB.scala 63:35]
  wire  _T_48 = valid_10 & _T_47; // @[TLB.scala 63:20]
  wire  _GEN_185 = _T_48 | _GEN_174; // @[TLB.scala 63:44]
  wire  _GEN_189 = _T_48 ? data_entry_r__T_49_data : _GEN_178; // @[TLB.scala 63:44]
  wire  _GEN_190 = _T_48 ? data_entry_w__T_49_data : _GEN_179; // @[TLB.scala 63:44]
  wire  _GEN_191 = _T_48 ? data_entry_x__T_49_data : _GEN_180; // @[TLB.scala 63:44]
  wire  _GEN_192 = _T_48 ? data_entry_u__T_49_data : _GEN_181; // @[TLB.scala 63:44]
  wire  _GEN_193 = _T_48 ? data_entry_a__T_49_data : _GEN_182; // @[TLB.scala 63:44]
  wire  _GEN_194 = _T_48 ? data_entry_d__T_49_data : _GEN_183; // @[TLB.scala 63:44]
  wire [21:0] _GEN_195 = _T_48 ? data_entry_ppn__T_49_data : _GEN_184; // @[TLB.scala 63:44]
  wire  _T_51 = data_vpn__T_50_data == vpn; // @[TLB.scala 63:35]
  wire  _T_52 = valid_11 & _T_51; // @[TLB.scala 63:20]
  wire  _GEN_196 = _T_52 | _GEN_185; // @[TLB.scala 63:44]
  wire  _GEN_200 = _T_52 ? data_entry_r__T_53_data : _GEN_189; // @[TLB.scala 63:44]
  wire  _GEN_201 = _T_52 ? data_entry_w__T_53_data : _GEN_190; // @[TLB.scala 63:44]
  wire  _GEN_202 = _T_52 ? data_entry_x__T_53_data : _GEN_191; // @[TLB.scala 63:44]
  wire  _GEN_203 = _T_52 ? data_entry_u__T_53_data : _GEN_192; // @[TLB.scala 63:44]
  wire  _GEN_204 = _T_52 ? data_entry_a__T_53_data : _GEN_193; // @[TLB.scala 63:44]
  wire  _GEN_205 = _T_52 ? data_entry_d__T_53_data : _GEN_194; // @[TLB.scala 63:44]
  wire [21:0] _GEN_206 = _T_52 ? data_entry_ppn__T_53_data : _GEN_195; // @[TLB.scala 63:44]
  wire  _T_55 = data_vpn__T_54_data == vpn; // @[TLB.scala 63:35]
  wire  _T_56 = valid_12 & _T_55; // @[TLB.scala 63:20]
  wire  _GEN_207 = _T_56 | _GEN_196; // @[TLB.scala 63:44]
  wire  _GEN_211 = _T_56 ? data_entry_r__T_57_data : _GEN_200; // @[TLB.scala 63:44]
  wire  _GEN_212 = _T_56 ? data_entry_w__T_57_data : _GEN_201; // @[TLB.scala 63:44]
  wire  _GEN_213 = _T_56 ? data_entry_x__T_57_data : _GEN_202; // @[TLB.scala 63:44]
  wire  _GEN_214 = _T_56 ? data_entry_u__T_57_data : _GEN_203; // @[TLB.scala 63:44]
  wire  _GEN_215 = _T_56 ? data_entry_a__T_57_data : _GEN_204; // @[TLB.scala 63:44]
  wire  _GEN_216 = _T_56 ? data_entry_d__T_57_data : _GEN_205; // @[TLB.scala 63:44]
  wire [21:0] _GEN_217 = _T_56 ? data_entry_ppn__T_57_data : _GEN_206; // @[TLB.scala 63:44]
  wire  _T_59 = data_vpn__T_58_data == vpn; // @[TLB.scala 63:35]
  wire  _T_60 = valid_13 & _T_59; // @[TLB.scala 63:20]
  wire  _GEN_218 = _T_60 | _GEN_207; // @[TLB.scala 63:44]
  wire  _GEN_222 = _T_60 ? data_entry_r__T_61_data : _GEN_211; // @[TLB.scala 63:44]
  wire  _GEN_223 = _T_60 ? data_entry_w__T_61_data : _GEN_212; // @[TLB.scala 63:44]
  wire  _GEN_224 = _T_60 ? data_entry_x__T_61_data : _GEN_213; // @[TLB.scala 63:44]
  wire  _GEN_225 = _T_60 ? data_entry_u__T_61_data : _GEN_214; // @[TLB.scala 63:44]
  wire  _GEN_226 = _T_60 ? data_entry_a__T_61_data : _GEN_215; // @[TLB.scala 63:44]
  wire  _GEN_227 = _T_60 ? data_entry_d__T_61_data : _GEN_216; // @[TLB.scala 63:44]
  wire [21:0] _GEN_228 = _T_60 ? data_entry_ppn__T_61_data : _GEN_217; // @[TLB.scala 63:44]
  wire  _T_63 = data_vpn__T_62_data == vpn; // @[TLB.scala 63:35]
  wire  _T_64 = valid_14 & _T_63; // @[TLB.scala 63:20]
  wire  _GEN_229 = _T_64 | _GEN_218; // @[TLB.scala 63:44]
  wire  _GEN_233 = _T_64 ? data_entry_r__T_65_data : _GEN_222; // @[TLB.scala 63:44]
  wire  _GEN_234 = _T_64 ? data_entry_w__T_65_data : _GEN_223; // @[TLB.scala 63:44]
  wire  _GEN_235 = _T_64 ? data_entry_x__T_65_data : _GEN_224; // @[TLB.scala 63:44]
  wire  _GEN_236 = _T_64 ? data_entry_u__T_65_data : _GEN_225; // @[TLB.scala 63:44]
  wire  _GEN_237 = _T_64 ? data_entry_a__T_65_data : _GEN_226; // @[TLB.scala 63:44]
  wire  _GEN_238 = _T_64 ? data_entry_d__T_65_data : _GEN_227; // @[TLB.scala 63:44]
  wire [21:0] _GEN_239 = _T_64 ? data_entry_ppn__T_65_data : _GEN_228; // @[TLB.scala 63:44]
  wire  _T_67 = data_vpn__T_66_data == vpn; // @[TLB.scala 63:35]
  wire  _T_68 = valid_15 & _T_67; // @[TLB.scala 63:20]
  assign data_vpn__T_6_addr = 4'h0;
  assign data_vpn__T_6_data = data_vpn[data_vpn__T_6_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_9_addr = 4'h0;
  assign data_vpn__T_9_data = data_vpn[data_vpn__T_9_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_10_addr = 4'h1;
  assign data_vpn__T_10_data = data_vpn[data_vpn__T_10_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_13_addr = 4'h1;
  assign data_vpn__T_13_data = data_vpn[data_vpn__T_13_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_14_addr = 4'h2;
  assign data_vpn__T_14_data = data_vpn[data_vpn__T_14_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_17_addr = 4'h2;
  assign data_vpn__T_17_data = data_vpn[data_vpn__T_17_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_18_addr = 4'h3;
  assign data_vpn__T_18_data = data_vpn[data_vpn__T_18_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_21_addr = 4'h3;
  assign data_vpn__T_21_data = data_vpn[data_vpn__T_21_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_22_addr = 4'h4;
  assign data_vpn__T_22_data = data_vpn[data_vpn__T_22_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_25_addr = 4'h4;
  assign data_vpn__T_25_data = data_vpn[data_vpn__T_25_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_26_addr = 4'h5;
  assign data_vpn__T_26_data = data_vpn[data_vpn__T_26_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_29_addr = 4'h5;
  assign data_vpn__T_29_data = data_vpn[data_vpn__T_29_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_30_addr = 4'h6;
  assign data_vpn__T_30_data = data_vpn[data_vpn__T_30_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_33_addr = 4'h6;
  assign data_vpn__T_33_data = data_vpn[data_vpn__T_33_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_34_addr = 4'h7;
  assign data_vpn__T_34_data = data_vpn[data_vpn__T_34_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_37_addr = 4'h7;
  assign data_vpn__T_37_data = data_vpn[data_vpn__T_37_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_38_addr = 4'h8;
  assign data_vpn__T_38_data = data_vpn[data_vpn__T_38_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_41_addr = 4'h8;
  assign data_vpn__T_41_data = data_vpn[data_vpn__T_41_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_42_addr = 4'h9;
  assign data_vpn__T_42_data = data_vpn[data_vpn__T_42_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_45_addr = 4'h9;
  assign data_vpn__T_45_data = data_vpn[data_vpn__T_45_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_46_addr = 4'ha;
  assign data_vpn__T_46_data = data_vpn[data_vpn__T_46_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_49_addr = 4'ha;
  assign data_vpn__T_49_data = data_vpn[data_vpn__T_49_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_50_addr = 4'hb;
  assign data_vpn__T_50_data = data_vpn[data_vpn__T_50_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_53_addr = 4'hb;
  assign data_vpn__T_53_data = data_vpn[data_vpn__T_53_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_54_addr = 4'hc;
  assign data_vpn__T_54_data = data_vpn[data_vpn__T_54_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_57_addr = 4'hc;
  assign data_vpn__T_57_data = data_vpn[data_vpn__T_57_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_58_addr = 4'hd;
  assign data_vpn__T_58_data = data_vpn[data_vpn__T_58_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_61_addr = 4'hd;
  assign data_vpn__T_61_data = data_vpn[data_vpn__T_61_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_62_addr = 4'he;
  assign data_vpn__T_62_data = data_vpn[data_vpn__T_62_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_65_addr = 4'he;
  assign data_vpn__T_65_data = data_vpn[data_vpn__T_65_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_66_addr = 4'hf;
  assign data_vpn__T_66_data = data_vpn[data_vpn__T_66_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_69_addr = 4'hf;
  assign data_vpn__T_69_data = data_vpn[data_vpn__T_69_addr]; // @[TLB.scala 37:18]
  assign data_vpn__T_1_data = io_vaddr[31:12];
  assign data_vpn__T_1_addr = pointer;
  assign data_vpn__T_1_mask = 1'h1;
  assign data_vpn__T_1_en = io_flush ? 1'h0 : io_wen;
  assign data_vpn__T_2_data = 20'h0;
  assign data_vpn__T_2_addr = pointer;
  assign data_vpn__T_2_mask = 1'h0;
  assign data_vpn__T_2_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_ppn__T_6_addr = 4'h0;
  assign data_entry_ppn__T_6_data = data_entry_ppn[data_entry_ppn__T_6_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_9_addr = 4'h0;
  assign data_entry_ppn__T_9_data = data_entry_ppn[data_entry_ppn__T_9_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_10_addr = 4'h1;
  assign data_entry_ppn__T_10_data = data_entry_ppn[data_entry_ppn__T_10_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_13_addr = 4'h1;
  assign data_entry_ppn__T_13_data = data_entry_ppn[data_entry_ppn__T_13_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_14_addr = 4'h2;
  assign data_entry_ppn__T_14_data = data_entry_ppn[data_entry_ppn__T_14_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_17_addr = 4'h2;
  assign data_entry_ppn__T_17_data = data_entry_ppn[data_entry_ppn__T_17_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_18_addr = 4'h3;
  assign data_entry_ppn__T_18_data = data_entry_ppn[data_entry_ppn__T_18_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_21_addr = 4'h3;
  assign data_entry_ppn__T_21_data = data_entry_ppn[data_entry_ppn__T_21_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_22_addr = 4'h4;
  assign data_entry_ppn__T_22_data = data_entry_ppn[data_entry_ppn__T_22_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_25_addr = 4'h4;
  assign data_entry_ppn__T_25_data = data_entry_ppn[data_entry_ppn__T_25_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_26_addr = 4'h5;
  assign data_entry_ppn__T_26_data = data_entry_ppn[data_entry_ppn__T_26_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_29_addr = 4'h5;
  assign data_entry_ppn__T_29_data = data_entry_ppn[data_entry_ppn__T_29_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_30_addr = 4'h6;
  assign data_entry_ppn__T_30_data = data_entry_ppn[data_entry_ppn__T_30_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_33_addr = 4'h6;
  assign data_entry_ppn__T_33_data = data_entry_ppn[data_entry_ppn__T_33_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_34_addr = 4'h7;
  assign data_entry_ppn__T_34_data = data_entry_ppn[data_entry_ppn__T_34_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_37_addr = 4'h7;
  assign data_entry_ppn__T_37_data = data_entry_ppn[data_entry_ppn__T_37_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_38_addr = 4'h8;
  assign data_entry_ppn__T_38_data = data_entry_ppn[data_entry_ppn__T_38_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_41_addr = 4'h8;
  assign data_entry_ppn__T_41_data = data_entry_ppn[data_entry_ppn__T_41_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_42_addr = 4'h9;
  assign data_entry_ppn__T_42_data = data_entry_ppn[data_entry_ppn__T_42_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_45_addr = 4'h9;
  assign data_entry_ppn__T_45_data = data_entry_ppn[data_entry_ppn__T_45_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_46_addr = 4'ha;
  assign data_entry_ppn__T_46_data = data_entry_ppn[data_entry_ppn__T_46_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_49_addr = 4'ha;
  assign data_entry_ppn__T_49_data = data_entry_ppn[data_entry_ppn__T_49_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_50_addr = 4'hb;
  assign data_entry_ppn__T_50_data = data_entry_ppn[data_entry_ppn__T_50_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_53_addr = 4'hb;
  assign data_entry_ppn__T_53_data = data_entry_ppn[data_entry_ppn__T_53_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_54_addr = 4'hc;
  assign data_entry_ppn__T_54_data = data_entry_ppn[data_entry_ppn__T_54_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_57_addr = 4'hc;
  assign data_entry_ppn__T_57_data = data_entry_ppn[data_entry_ppn__T_57_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_58_addr = 4'hd;
  assign data_entry_ppn__T_58_data = data_entry_ppn[data_entry_ppn__T_58_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_61_addr = 4'hd;
  assign data_entry_ppn__T_61_data = data_entry_ppn[data_entry_ppn__T_61_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_62_addr = 4'he;
  assign data_entry_ppn__T_62_data = data_entry_ppn[data_entry_ppn__T_62_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_65_addr = 4'he;
  assign data_entry_ppn__T_65_data = data_entry_ppn[data_entry_ppn__T_65_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_66_addr = 4'hf;
  assign data_entry_ppn__T_66_data = data_entry_ppn[data_entry_ppn__T_66_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_69_addr = 4'hf;
  assign data_entry_ppn__T_69_data = data_entry_ppn[data_entry_ppn__T_69_addr]; // @[TLB.scala 37:18]
  assign data_entry_ppn__T_1_data = 22'h0;
  assign data_entry_ppn__T_1_addr = pointer;
  assign data_entry_ppn__T_1_mask = 1'h0;
  assign data_entry_ppn__T_1_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_ppn__T_2_data = io_went_ppn;
  assign data_entry_ppn__T_2_addr = pointer;
  assign data_entry_ppn__T_2_mask = 1'h1;
  assign data_entry_ppn__T_2_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_d__T_6_addr = 4'h0;
  assign data_entry_d__T_6_data = data_entry_d[data_entry_d__T_6_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_9_addr = 4'h0;
  assign data_entry_d__T_9_data = data_entry_d[data_entry_d__T_9_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_10_addr = 4'h1;
  assign data_entry_d__T_10_data = data_entry_d[data_entry_d__T_10_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_13_addr = 4'h1;
  assign data_entry_d__T_13_data = data_entry_d[data_entry_d__T_13_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_14_addr = 4'h2;
  assign data_entry_d__T_14_data = data_entry_d[data_entry_d__T_14_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_17_addr = 4'h2;
  assign data_entry_d__T_17_data = data_entry_d[data_entry_d__T_17_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_18_addr = 4'h3;
  assign data_entry_d__T_18_data = data_entry_d[data_entry_d__T_18_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_21_addr = 4'h3;
  assign data_entry_d__T_21_data = data_entry_d[data_entry_d__T_21_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_22_addr = 4'h4;
  assign data_entry_d__T_22_data = data_entry_d[data_entry_d__T_22_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_25_addr = 4'h4;
  assign data_entry_d__T_25_data = data_entry_d[data_entry_d__T_25_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_26_addr = 4'h5;
  assign data_entry_d__T_26_data = data_entry_d[data_entry_d__T_26_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_29_addr = 4'h5;
  assign data_entry_d__T_29_data = data_entry_d[data_entry_d__T_29_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_30_addr = 4'h6;
  assign data_entry_d__T_30_data = data_entry_d[data_entry_d__T_30_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_33_addr = 4'h6;
  assign data_entry_d__T_33_data = data_entry_d[data_entry_d__T_33_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_34_addr = 4'h7;
  assign data_entry_d__T_34_data = data_entry_d[data_entry_d__T_34_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_37_addr = 4'h7;
  assign data_entry_d__T_37_data = data_entry_d[data_entry_d__T_37_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_38_addr = 4'h8;
  assign data_entry_d__T_38_data = data_entry_d[data_entry_d__T_38_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_41_addr = 4'h8;
  assign data_entry_d__T_41_data = data_entry_d[data_entry_d__T_41_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_42_addr = 4'h9;
  assign data_entry_d__T_42_data = data_entry_d[data_entry_d__T_42_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_45_addr = 4'h9;
  assign data_entry_d__T_45_data = data_entry_d[data_entry_d__T_45_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_46_addr = 4'ha;
  assign data_entry_d__T_46_data = data_entry_d[data_entry_d__T_46_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_49_addr = 4'ha;
  assign data_entry_d__T_49_data = data_entry_d[data_entry_d__T_49_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_50_addr = 4'hb;
  assign data_entry_d__T_50_data = data_entry_d[data_entry_d__T_50_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_53_addr = 4'hb;
  assign data_entry_d__T_53_data = data_entry_d[data_entry_d__T_53_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_54_addr = 4'hc;
  assign data_entry_d__T_54_data = data_entry_d[data_entry_d__T_54_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_57_addr = 4'hc;
  assign data_entry_d__T_57_data = data_entry_d[data_entry_d__T_57_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_58_addr = 4'hd;
  assign data_entry_d__T_58_data = data_entry_d[data_entry_d__T_58_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_61_addr = 4'hd;
  assign data_entry_d__T_61_data = data_entry_d[data_entry_d__T_61_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_62_addr = 4'he;
  assign data_entry_d__T_62_data = data_entry_d[data_entry_d__T_62_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_65_addr = 4'he;
  assign data_entry_d__T_65_data = data_entry_d[data_entry_d__T_65_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_66_addr = 4'hf;
  assign data_entry_d__T_66_data = data_entry_d[data_entry_d__T_66_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_69_addr = 4'hf;
  assign data_entry_d__T_69_data = data_entry_d[data_entry_d__T_69_addr]; // @[TLB.scala 37:18]
  assign data_entry_d__T_1_data = 1'h0;
  assign data_entry_d__T_1_addr = pointer;
  assign data_entry_d__T_1_mask = 1'h0;
  assign data_entry_d__T_1_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_d__T_2_data = io_went_d;
  assign data_entry_d__T_2_addr = pointer;
  assign data_entry_d__T_2_mask = 1'h1;
  assign data_entry_d__T_2_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_a__T_6_addr = 4'h0;
  assign data_entry_a__T_6_data = data_entry_a[data_entry_a__T_6_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_9_addr = 4'h0;
  assign data_entry_a__T_9_data = data_entry_a[data_entry_a__T_9_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_10_addr = 4'h1;
  assign data_entry_a__T_10_data = data_entry_a[data_entry_a__T_10_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_13_addr = 4'h1;
  assign data_entry_a__T_13_data = data_entry_a[data_entry_a__T_13_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_14_addr = 4'h2;
  assign data_entry_a__T_14_data = data_entry_a[data_entry_a__T_14_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_17_addr = 4'h2;
  assign data_entry_a__T_17_data = data_entry_a[data_entry_a__T_17_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_18_addr = 4'h3;
  assign data_entry_a__T_18_data = data_entry_a[data_entry_a__T_18_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_21_addr = 4'h3;
  assign data_entry_a__T_21_data = data_entry_a[data_entry_a__T_21_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_22_addr = 4'h4;
  assign data_entry_a__T_22_data = data_entry_a[data_entry_a__T_22_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_25_addr = 4'h4;
  assign data_entry_a__T_25_data = data_entry_a[data_entry_a__T_25_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_26_addr = 4'h5;
  assign data_entry_a__T_26_data = data_entry_a[data_entry_a__T_26_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_29_addr = 4'h5;
  assign data_entry_a__T_29_data = data_entry_a[data_entry_a__T_29_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_30_addr = 4'h6;
  assign data_entry_a__T_30_data = data_entry_a[data_entry_a__T_30_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_33_addr = 4'h6;
  assign data_entry_a__T_33_data = data_entry_a[data_entry_a__T_33_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_34_addr = 4'h7;
  assign data_entry_a__T_34_data = data_entry_a[data_entry_a__T_34_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_37_addr = 4'h7;
  assign data_entry_a__T_37_data = data_entry_a[data_entry_a__T_37_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_38_addr = 4'h8;
  assign data_entry_a__T_38_data = data_entry_a[data_entry_a__T_38_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_41_addr = 4'h8;
  assign data_entry_a__T_41_data = data_entry_a[data_entry_a__T_41_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_42_addr = 4'h9;
  assign data_entry_a__T_42_data = data_entry_a[data_entry_a__T_42_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_45_addr = 4'h9;
  assign data_entry_a__T_45_data = data_entry_a[data_entry_a__T_45_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_46_addr = 4'ha;
  assign data_entry_a__T_46_data = data_entry_a[data_entry_a__T_46_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_49_addr = 4'ha;
  assign data_entry_a__T_49_data = data_entry_a[data_entry_a__T_49_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_50_addr = 4'hb;
  assign data_entry_a__T_50_data = data_entry_a[data_entry_a__T_50_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_53_addr = 4'hb;
  assign data_entry_a__T_53_data = data_entry_a[data_entry_a__T_53_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_54_addr = 4'hc;
  assign data_entry_a__T_54_data = data_entry_a[data_entry_a__T_54_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_57_addr = 4'hc;
  assign data_entry_a__T_57_data = data_entry_a[data_entry_a__T_57_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_58_addr = 4'hd;
  assign data_entry_a__T_58_data = data_entry_a[data_entry_a__T_58_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_61_addr = 4'hd;
  assign data_entry_a__T_61_data = data_entry_a[data_entry_a__T_61_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_62_addr = 4'he;
  assign data_entry_a__T_62_data = data_entry_a[data_entry_a__T_62_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_65_addr = 4'he;
  assign data_entry_a__T_65_data = data_entry_a[data_entry_a__T_65_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_66_addr = 4'hf;
  assign data_entry_a__T_66_data = data_entry_a[data_entry_a__T_66_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_69_addr = 4'hf;
  assign data_entry_a__T_69_data = data_entry_a[data_entry_a__T_69_addr]; // @[TLB.scala 37:18]
  assign data_entry_a__T_1_data = 1'h0;
  assign data_entry_a__T_1_addr = pointer;
  assign data_entry_a__T_1_mask = 1'h0;
  assign data_entry_a__T_1_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_a__T_2_data = io_went_a;
  assign data_entry_a__T_2_addr = pointer;
  assign data_entry_a__T_2_mask = 1'h1;
  assign data_entry_a__T_2_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_u__T_6_addr = 4'h0;
  assign data_entry_u__T_6_data = data_entry_u[data_entry_u__T_6_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_9_addr = 4'h0;
  assign data_entry_u__T_9_data = data_entry_u[data_entry_u__T_9_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_10_addr = 4'h1;
  assign data_entry_u__T_10_data = data_entry_u[data_entry_u__T_10_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_13_addr = 4'h1;
  assign data_entry_u__T_13_data = data_entry_u[data_entry_u__T_13_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_14_addr = 4'h2;
  assign data_entry_u__T_14_data = data_entry_u[data_entry_u__T_14_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_17_addr = 4'h2;
  assign data_entry_u__T_17_data = data_entry_u[data_entry_u__T_17_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_18_addr = 4'h3;
  assign data_entry_u__T_18_data = data_entry_u[data_entry_u__T_18_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_21_addr = 4'h3;
  assign data_entry_u__T_21_data = data_entry_u[data_entry_u__T_21_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_22_addr = 4'h4;
  assign data_entry_u__T_22_data = data_entry_u[data_entry_u__T_22_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_25_addr = 4'h4;
  assign data_entry_u__T_25_data = data_entry_u[data_entry_u__T_25_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_26_addr = 4'h5;
  assign data_entry_u__T_26_data = data_entry_u[data_entry_u__T_26_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_29_addr = 4'h5;
  assign data_entry_u__T_29_data = data_entry_u[data_entry_u__T_29_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_30_addr = 4'h6;
  assign data_entry_u__T_30_data = data_entry_u[data_entry_u__T_30_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_33_addr = 4'h6;
  assign data_entry_u__T_33_data = data_entry_u[data_entry_u__T_33_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_34_addr = 4'h7;
  assign data_entry_u__T_34_data = data_entry_u[data_entry_u__T_34_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_37_addr = 4'h7;
  assign data_entry_u__T_37_data = data_entry_u[data_entry_u__T_37_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_38_addr = 4'h8;
  assign data_entry_u__T_38_data = data_entry_u[data_entry_u__T_38_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_41_addr = 4'h8;
  assign data_entry_u__T_41_data = data_entry_u[data_entry_u__T_41_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_42_addr = 4'h9;
  assign data_entry_u__T_42_data = data_entry_u[data_entry_u__T_42_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_45_addr = 4'h9;
  assign data_entry_u__T_45_data = data_entry_u[data_entry_u__T_45_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_46_addr = 4'ha;
  assign data_entry_u__T_46_data = data_entry_u[data_entry_u__T_46_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_49_addr = 4'ha;
  assign data_entry_u__T_49_data = data_entry_u[data_entry_u__T_49_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_50_addr = 4'hb;
  assign data_entry_u__T_50_data = data_entry_u[data_entry_u__T_50_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_53_addr = 4'hb;
  assign data_entry_u__T_53_data = data_entry_u[data_entry_u__T_53_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_54_addr = 4'hc;
  assign data_entry_u__T_54_data = data_entry_u[data_entry_u__T_54_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_57_addr = 4'hc;
  assign data_entry_u__T_57_data = data_entry_u[data_entry_u__T_57_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_58_addr = 4'hd;
  assign data_entry_u__T_58_data = data_entry_u[data_entry_u__T_58_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_61_addr = 4'hd;
  assign data_entry_u__T_61_data = data_entry_u[data_entry_u__T_61_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_62_addr = 4'he;
  assign data_entry_u__T_62_data = data_entry_u[data_entry_u__T_62_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_65_addr = 4'he;
  assign data_entry_u__T_65_data = data_entry_u[data_entry_u__T_65_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_66_addr = 4'hf;
  assign data_entry_u__T_66_data = data_entry_u[data_entry_u__T_66_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_69_addr = 4'hf;
  assign data_entry_u__T_69_data = data_entry_u[data_entry_u__T_69_addr]; // @[TLB.scala 37:18]
  assign data_entry_u__T_1_data = 1'h0;
  assign data_entry_u__T_1_addr = pointer;
  assign data_entry_u__T_1_mask = 1'h0;
  assign data_entry_u__T_1_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_u__T_2_data = io_went_u;
  assign data_entry_u__T_2_addr = pointer;
  assign data_entry_u__T_2_mask = 1'h1;
  assign data_entry_u__T_2_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_x__T_6_addr = 4'h0;
  assign data_entry_x__T_6_data = data_entry_x[data_entry_x__T_6_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_9_addr = 4'h0;
  assign data_entry_x__T_9_data = data_entry_x[data_entry_x__T_9_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_10_addr = 4'h1;
  assign data_entry_x__T_10_data = data_entry_x[data_entry_x__T_10_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_13_addr = 4'h1;
  assign data_entry_x__T_13_data = data_entry_x[data_entry_x__T_13_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_14_addr = 4'h2;
  assign data_entry_x__T_14_data = data_entry_x[data_entry_x__T_14_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_17_addr = 4'h2;
  assign data_entry_x__T_17_data = data_entry_x[data_entry_x__T_17_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_18_addr = 4'h3;
  assign data_entry_x__T_18_data = data_entry_x[data_entry_x__T_18_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_21_addr = 4'h3;
  assign data_entry_x__T_21_data = data_entry_x[data_entry_x__T_21_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_22_addr = 4'h4;
  assign data_entry_x__T_22_data = data_entry_x[data_entry_x__T_22_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_25_addr = 4'h4;
  assign data_entry_x__T_25_data = data_entry_x[data_entry_x__T_25_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_26_addr = 4'h5;
  assign data_entry_x__T_26_data = data_entry_x[data_entry_x__T_26_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_29_addr = 4'h5;
  assign data_entry_x__T_29_data = data_entry_x[data_entry_x__T_29_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_30_addr = 4'h6;
  assign data_entry_x__T_30_data = data_entry_x[data_entry_x__T_30_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_33_addr = 4'h6;
  assign data_entry_x__T_33_data = data_entry_x[data_entry_x__T_33_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_34_addr = 4'h7;
  assign data_entry_x__T_34_data = data_entry_x[data_entry_x__T_34_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_37_addr = 4'h7;
  assign data_entry_x__T_37_data = data_entry_x[data_entry_x__T_37_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_38_addr = 4'h8;
  assign data_entry_x__T_38_data = data_entry_x[data_entry_x__T_38_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_41_addr = 4'h8;
  assign data_entry_x__T_41_data = data_entry_x[data_entry_x__T_41_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_42_addr = 4'h9;
  assign data_entry_x__T_42_data = data_entry_x[data_entry_x__T_42_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_45_addr = 4'h9;
  assign data_entry_x__T_45_data = data_entry_x[data_entry_x__T_45_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_46_addr = 4'ha;
  assign data_entry_x__T_46_data = data_entry_x[data_entry_x__T_46_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_49_addr = 4'ha;
  assign data_entry_x__T_49_data = data_entry_x[data_entry_x__T_49_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_50_addr = 4'hb;
  assign data_entry_x__T_50_data = data_entry_x[data_entry_x__T_50_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_53_addr = 4'hb;
  assign data_entry_x__T_53_data = data_entry_x[data_entry_x__T_53_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_54_addr = 4'hc;
  assign data_entry_x__T_54_data = data_entry_x[data_entry_x__T_54_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_57_addr = 4'hc;
  assign data_entry_x__T_57_data = data_entry_x[data_entry_x__T_57_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_58_addr = 4'hd;
  assign data_entry_x__T_58_data = data_entry_x[data_entry_x__T_58_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_61_addr = 4'hd;
  assign data_entry_x__T_61_data = data_entry_x[data_entry_x__T_61_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_62_addr = 4'he;
  assign data_entry_x__T_62_data = data_entry_x[data_entry_x__T_62_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_65_addr = 4'he;
  assign data_entry_x__T_65_data = data_entry_x[data_entry_x__T_65_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_66_addr = 4'hf;
  assign data_entry_x__T_66_data = data_entry_x[data_entry_x__T_66_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_69_addr = 4'hf;
  assign data_entry_x__T_69_data = data_entry_x[data_entry_x__T_69_addr]; // @[TLB.scala 37:18]
  assign data_entry_x__T_1_data = 1'h0;
  assign data_entry_x__T_1_addr = pointer;
  assign data_entry_x__T_1_mask = 1'h0;
  assign data_entry_x__T_1_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_x__T_2_data = io_went_x;
  assign data_entry_x__T_2_addr = pointer;
  assign data_entry_x__T_2_mask = 1'h1;
  assign data_entry_x__T_2_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_w__T_6_addr = 4'h0;
  assign data_entry_w__T_6_data = data_entry_w[data_entry_w__T_6_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_9_addr = 4'h0;
  assign data_entry_w__T_9_data = data_entry_w[data_entry_w__T_9_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_10_addr = 4'h1;
  assign data_entry_w__T_10_data = data_entry_w[data_entry_w__T_10_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_13_addr = 4'h1;
  assign data_entry_w__T_13_data = data_entry_w[data_entry_w__T_13_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_14_addr = 4'h2;
  assign data_entry_w__T_14_data = data_entry_w[data_entry_w__T_14_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_17_addr = 4'h2;
  assign data_entry_w__T_17_data = data_entry_w[data_entry_w__T_17_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_18_addr = 4'h3;
  assign data_entry_w__T_18_data = data_entry_w[data_entry_w__T_18_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_21_addr = 4'h3;
  assign data_entry_w__T_21_data = data_entry_w[data_entry_w__T_21_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_22_addr = 4'h4;
  assign data_entry_w__T_22_data = data_entry_w[data_entry_w__T_22_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_25_addr = 4'h4;
  assign data_entry_w__T_25_data = data_entry_w[data_entry_w__T_25_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_26_addr = 4'h5;
  assign data_entry_w__T_26_data = data_entry_w[data_entry_w__T_26_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_29_addr = 4'h5;
  assign data_entry_w__T_29_data = data_entry_w[data_entry_w__T_29_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_30_addr = 4'h6;
  assign data_entry_w__T_30_data = data_entry_w[data_entry_w__T_30_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_33_addr = 4'h6;
  assign data_entry_w__T_33_data = data_entry_w[data_entry_w__T_33_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_34_addr = 4'h7;
  assign data_entry_w__T_34_data = data_entry_w[data_entry_w__T_34_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_37_addr = 4'h7;
  assign data_entry_w__T_37_data = data_entry_w[data_entry_w__T_37_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_38_addr = 4'h8;
  assign data_entry_w__T_38_data = data_entry_w[data_entry_w__T_38_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_41_addr = 4'h8;
  assign data_entry_w__T_41_data = data_entry_w[data_entry_w__T_41_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_42_addr = 4'h9;
  assign data_entry_w__T_42_data = data_entry_w[data_entry_w__T_42_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_45_addr = 4'h9;
  assign data_entry_w__T_45_data = data_entry_w[data_entry_w__T_45_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_46_addr = 4'ha;
  assign data_entry_w__T_46_data = data_entry_w[data_entry_w__T_46_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_49_addr = 4'ha;
  assign data_entry_w__T_49_data = data_entry_w[data_entry_w__T_49_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_50_addr = 4'hb;
  assign data_entry_w__T_50_data = data_entry_w[data_entry_w__T_50_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_53_addr = 4'hb;
  assign data_entry_w__T_53_data = data_entry_w[data_entry_w__T_53_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_54_addr = 4'hc;
  assign data_entry_w__T_54_data = data_entry_w[data_entry_w__T_54_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_57_addr = 4'hc;
  assign data_entry_w__T_57_data = data_entry_w[data_entry_w__T_57_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_58_addr = 4'hd;
  assign data_entry_w__T_58_data = data_entry_w[data_entry_w__T_58_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_61_addr = 4'hd;
  assign data_entry_w__T_61_data = data_entry_w[data_entry_w__T_61_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_62_addr = 4'he;
  assign data_entry_w__T_62_data = data_entry_w[data_entry_w__T_62_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_65_addr = 4'he;
  assign data_entry_w__T_65_data = data_entry_w[data_entry_w__T_65_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_66_addr = 4'hf;
  assign data_entry_w__T_66_data = data_entry_w[data_entry_w__T_66_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_69_addr = 4'hf;
  assign data_entry_w__T_69_data = data_entry_w[data_entry_w__T_69_addr]; // @[TLB.scala 37:18]
  assign data_entry_w__T_1_data = 1'h0;
  assign data_entry_w__T_1_addr = pointer;
  assign data_entry_w__T_1_mask = 1'h0;
  assign data_entry_w__T_1_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_w__T_2_data = io_went_w;
  assign data_entry_w__T_2_addr = pointer;
  assign data_entry_w__T_2_mask = 1'h1;
  assign data_entry_w__T_2_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_r__T_6_addr = 4'h0;
  assign data_entry_r__T_6_data = data_entry_r[data_entry_r__T_6_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_9_addr = 4'h0;
  assign data_entry_r__T_9_data = data_entry_r[data_entry_r__T_9_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_10_addr = 4'h1;
  assign data_entry_r__T_10_data = data_entry_r[data_entry_r__T_10_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_13_addr = 4'h1;
  assign data_entry_r__T_13_data = data_entry_r[data_entry_r__T_13_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_14_addr = 4'h2;
  assign data_entry_r__T_14_data = data_entry_r[data_entry_r__T_14_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_17_addr = 4'h2;
  assign data_entry_r__T_17_data = data_entry_r[data_entry_r__T_17_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_18_addr = 4'h3;
  assign data_entry_r__T_18_data = data_entry_r[data_entry_r__T_18_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_21_addr = 4'h3;
  assign data_entry_r__T_21_data = data_entry_r[data_entry_r__T_21_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_22_addr = 4'h4;
  assign data_entry_r__T_22_data = data_entry_r[data_entry_r__T_22_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_25_addr = 4'h4;
  assign data_entry_r__T_25_data = data_entry_r[data_entry_r__T_25_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_26_addr = 4'h5;
  assign data_entry_r__T_26_data = data_entry_r[data_entry_r__T_26_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_29_addr = 4'h5;
  assign data_entry_r__T_29_data = data_entry_r[data_entry_r__T_29_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_30_addr = 4'h6;
  assign data_entry_r__T_30_data = data_entry_r[data_entry_r__T_30_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_33_addr = 4'h6;
  assign data_entry_r__T_33_data = data_entry_r[data_entry_r__T_33_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_34_addr = 4'h7;
  assign data_entry_r__T_34_data = data_entry_r[data_entry_r__T_34_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_37_addr = 4'h7;
  assign data_entry_r__T_37_data = data_entry_r[data_entry_r__T_37_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_38_addr = 4'h8;
  assign data_entry_r__T_38_data = data_entry_r[data_entry_r__T_38_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_41_addr = 4'h8;
  assign data_entry_r__T_41_data = data_entry_r[data_entry_r__T_41_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_42_addr = 4'h9;
  assign data_entry_r__T_42_data = data_entry_r[data_entry_r__T_42_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_45_addr = 4'h9;
  assign data_entry_r__T_45_data = data_entry_r[data_entry_r__T_45_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_46_addr = 4'ha;
  assign data_entry_r__T_46_data = data_entry_r[data_entry_r__T_46_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_49_addr = 4'ha;
  assign data_entry_r__T_49_data = data_entry_r[data_entry_r__T_49_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_50_addr = 4'hb;
  assign data_entry_r__T_50_data = data_entry_r[data_entry_r__T_50_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_53_addr = 4'hb;
  assign data_entry_r__T_53_data = data_entry_r[data_entry_r__T_53_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_54_addr = 4'hc;
  assign data_entry_r__T_54_data = data_entry_r[data_entry_r__T_54_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_57_addr = 4'hc;
  assign data_entry_r__T_57_data = data_entry_r[data_entry_r__T_57_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_58_addr = 4'hd;
  assign data_entry_r__T_58_data = data_entry_r[data_entry_r__T_58_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_61_addr = 4'hd;
  assign data_entry_r__T_61_data = data_entry_r[data_entry_r__T_61_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_62_addr = 4'he;
  assign data_entry_r__T_62_data = data_entry_r[data_entry_r__T_62_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_65_addr = 4'he;
  assign data_entry_r__T_65_data = data_entry_r[data_entry_r__T_65_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_66_addr = 4'hf;
  assign data_entry_r__T_66_data = data_entry_r[data_entry_r__T_66_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_69_addr = 4'hf;
  assign data_entry_r__T_69_data = data_entry_r[data_entry_r__T_69_addr]; // @[TLB.scala 37:18]
  assign data_entry_r__T_1_data = 1'h0;
  assign data_entry_r__T_1_addr = pointer;
  assign data_entry_r__T_1_mask = 1'h0;
  assign data_entry_r__T_1_en = io_flush ? 1'h0 : io_wen;
  assign data_entry_r__T_2_data = io_went_r;
  assign data_entry_r__T_2_addr = pointer;
  assign data_entry_r__T_2_mask = 1'h1;
  assign data_entry_r__T_2_en = io_flush ? 1'h0 : io_wen;
  assign io_valid = _T_68 | _GEN_229; // @[TLB.scala 70:13]
  assign io_rent_ppn = _T_68 ? data_entry_ppn__T_69_data : _GEN_239; // @[TLB.scala 71:13]
  assign io_rent_d = _T_68 ? data_entry_d__T_69_data : _GEN_238; // @[TLB.scala 71:13]
  assign io_rent_a = _T_68 ? data_entry_a__T_69_data : _GEN_237; // @[TLB.scala 71:13]
  assign io_rent_u = _T_68 ? data_entry_u__T_69_data : _GEN_236; // @[TLB.scala 71:13]
  assign io_rent_x = _T_68 ? data_entry_x__T_69_data : _GEN_235; // @[TLB.scala 71:13]
  assign io_rent_w = _T_68 ? data_entry_w__T_69_data : _GEN_234; // @[TLB.scala 71:13]
  assign io_rent_r = _T_68 ? data_entry_r__T_69_data : _GEN_233; // @[TLB.scala 71:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    data_vpn[initvar] = _RAND_0[19:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    data_entry_ppn[initvar] = _RAND_1[21:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_2 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    data_entry_d[initvar] = _RAND_2[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    data_entry_a[initvar] = _RAND_3[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_4 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    data_entry_u[initvar] = _RAND_4[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_5 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    data_entry_x[initvar] = _RAND_5[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    data_entry_w[initvar] = _RAND_6[0:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_7 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    data_entry_r[initvar] = _RAND_7[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  valid_0 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  valid_1 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  valid_2 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  valid_3 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  valid_4 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  valid_5 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  valid_6 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  valid_7 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  valid_8 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  valid_9 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  valid_10 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  valid_11 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valid_12 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  valid_13 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  valid_14 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  valid_15 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  pointer = _RAND_24[3:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(data_vpn__T_1_en & data_vpn__T_1_mask) begin
      data_vpn[data_vpn__T_1_addr] <= data_vpn__T_1_data; // @[TLB.scala 37:18]
    end
    if(data_vpn__T_2_en & data_vpn__T_2_mask) begin
      data_vpn[data_vpn__T_2_addr] <= data_vpn__T_2_data; // @[TLB.scala 37:18]
    end
    if(data_entry_ppn__T_1_en & data_entry_ppn__T_1_mask) begin
      data_entry_ppn[data_entry_ppn__T_1_addr] <= data_entry_ppn__T_1_data; // @[TLB.scala 37:18]
    end
    if(data_entry_ppn__T_2_en & data_entry_ppn__T_2_mask) begin
      data_entry_ppn[data_entry_ppn__T_2_addr] <= data_entry_ppn__T_2_data; // @[TLB.scala 37:18]
    end
    if(data_entry_d__T_1_en & data_entry_d__T_1_mask) begin
      data_entry_d[data_entry_d__T_1_addr] <= data_entry_d__T_1_data; // @[TLB.scala 37:18]
    end
    if(data_entry_d__T_2_en & data_entry_d__T_2_mask) begin
      data_entry_d[data_entry_d__T_2_addr] <= data_entry_d__T_2_data; // @[TLB.scala 37:18]
    end
    if(data_entry_a__T_1_en & data_entry_a__T_1_mask) begin
      data_entry_a[data_entry_a__T_1_addr] <= data_entry_a__T_1_data; // @[TLB.scala 37:18]
    end
    if(data_entry_a__T_2_en & data_entry_a__T_2_mask) begin
      data_entry_a[data_entry_a__T_2_addr] <= data_entry_a__T_2_data; // @[TLB.scala 37:18]
    end
    if(data_entry_u__T_1_en & data_entry_u__T_1_mask) begin
      data_entry_u[data_entry_u__T_1_addr] <= data_entry_u__T_1_data; // @[TLB.scala 37:18]
    end
    if(data_entry_u__T_2_en & data_entry_u__T_2_mask) begin
      data_entry_u[data_entry_u__T_2_addr] <= data_entry_u__T_2_data; // @[TLB.scala 37:18]
    end
    if(data_entry_x__T_1_en & data_entry_x__T_1_mask) begin
      data_entry_x[data_entry_x__T_1_addr] <= data_entry_x__T_1_data; // @[TLB.scala 37:18]
    end
    if(data_entry_x__T_2_en & data_entry_x__T_2_mask) begin
      data_entry_x[data_entry_x__T_2_addr] <= data_entry_x__T_2_data; // @[TLB.scala 37:18]
    end
    if(data_entry_w__T_1_en & data_entry_w__T_1_mask) begin
      data_entry_w[data_entry_w__T_1_addr] <= data_entry_w__T_1_data; // @[TLB.scala 37:18]
    end
    if(data_entry_w__T_2_en & data_entry_w__T_2_mask) begin
      data_entry_w[data_entry_w__T_2_addr] <= data_entry_w__T_2_data; // @[TLB.scala 37:18]
    end
    if(data_entry_r__T_1_en & data_entry_r__T_1_mask) begin
      data_entry_r[data_entry_r__T_1_addr] <= data_entry_r__T_1_data; // @[TLB.scala 37:18]
    end
    if(data_entry_r__T_2_en & data_entry_r__T_2_mask) begin
      data_entry_r[data_entry_r__T_2_addr] <= data_entry_r__T_2_data; // @[TLB.scala 37:18]
    end
    if (reset) begin
      valid_0 <= 1'h0;
    end else if (io_flush) begin
      valid_0 <= 1'h0;
    end else if (io_wen) begin
      valid_0 <= _GEN_0;
    end
    if (reset) begin
      valid_1 <= 1'h0;
    end else if (io_flush) begin
      valid_1 <= 1'h0;
    end else if (io_wen) begin
      valid_1 <= _GEN_1;
    end
    if (reset) begin
      valid_2 <= 1'h0;
    end else if (io_flush) begin
      valid_2 <= 1'h0;
    end else if (io_wen) begin
      valid_2 <= _GEN_2;
    end
    if (reset) begin
      valid_3 <= 1'h0;
    end else if (io_flush) begin
      valid_3 <= 1'h0;
    end else if (io_wen) begin
      valid_3 <= _GEN_3;
    end
    if (reset) begin
      valid_4 <= 1'h0;
    end else if (io_flush) begin
      valid_4 <= 1'h0;
    end else if (io_wen) begin
      valid_4 <= _GEN_4;
    end
    if (reset) begin
      valid_5 <= 1'h0;
    end else if (io_flush) begin
      valid_5 <= 1'h0;
    end else if (io_wen) begin
      valid_5 <= _GEN_5;
    end
    if (reset) begin
      valid_6 <= 1'h0;
    end else if (io_flush) begin
      valid_6 <= 1'h0;
    end else if (io_wen) begin
      valid_6 <= _GEN_6;
    end
    if (reset) begin
      valid_7 <= 1'h0;
    end else if (io_flush) begin
      valid_7 <= 1'h0;
    end else if (io_wen) begin
      valid_7 <= _GEN_7;
    end
    if (reset) begin
      valid_8 <= 1'h0;
    end else if (io_flush) begin
      valid_8 <= 1'h0;
    end else if (io_wen) begin
      valid_8 <= _GEN_8;
    end
    if (reset) begin
      valid_9 <= 1'h0;
    end else if (io_flush) begin
      valid_9 <= 1'h0;
    end else if (io_wen) begin
      valid_9 <= _GEN_9;
    end
    if (reset) begin
      valid_10 <= 1'h0;
    end else if (io_flush) begin
      valid_10 <= 1'h0;
    end else if (io_wen) begin
      valid_10 <= _GEN_10;
    end
    if (reset) begin
      valid_11 <= 1'h0;
    end else if (io_flush) begin
      valid_11 <= 1'h0;
    end else if (io_wen) begin
      valid_11 <= _GEN_11;
    end
    if (reset) begin
      valid_12 <= 1'h0;
    end else if (io_flush) begin
      valid_12 <= 1'h0;
    end else if (io_wen) begin
      valid_12 <= _GEN_12;
    end
    if (reset) begin
      valid_13 <= 1'h0;
    end else if (io_flush) begin
      valid_13 <= 1'h0;
    end else if (io_wen) begin
      valid_13 <= _GEN_13;
    end
    if (reset) begin
      valid_14 <= 1'h0;
    end else if (io_flush) begin
      valid_14 <= 1'h0;
    end else if (io_wen) begin
      valid_14 <= _GEN_14;
    end
    if (reset) begin
      valid_15 <= 1'h0;
    end else if (io_flush) begin
      valid_15 <= 1'h0;
    end else if (io_wen) begin
      valid_15 <= _GEN_15;
    end
    if (reset) begin
      pointer <= 4'h0;
    end else if (!(io_flush)) begin
      if (io_wen) begin
        pointer <= _T_4;
      end
    end
  end
endmodule
module MMU(
  input         clock,
  input         reset,
  input         io_en,
  input         io_flush,
  input  [21:0] io_basePpn,
  input         io_sum,
  input         io_smode,
  input  [31:0] io_vaddr,
  output        io_valid,
  output        io_fault,
  output [31:0] io_paddr,
  output        io_data_en,
  input         io_data_valid,
  output [31:0] io_data_addr,
  input  [31:0] io_data_rdata
);
  wire  tlb_clock; // @[MMU.scala 65:19]
  wire  tlb_reset; // @[MMU.scala 65:19]
  wire  tlb_io_flush; // @[MMU.scala 65:19]
  wire  tlb_io_wen; // @[MMU.scala 65:19]
  wire [31:0] tlb_io_vaddr; // @[MMU.scala 65:19]
  wire [21:0] tlb_io_went_ppn; // @[MMU.scala 65:19]
  wire  tlb_io_went_d; // @[MMU.scala 65:19]
  wire  tlb_io_went_a; // @[MMU.scala 65:19]
  wire  tlb_io_went_u; // @[MMU.scala 65:19]
  wire  tlb_io_went_x; // @[MMU.scala 65:19]
  wire  tlb_io_went_w; // @[MMU.scala 65:19]
  wire  tlb_io_went_r; // @[MMU.scala 65:19]
  wire  tlb_io_valid; // @[MMU.scala 65:19]
  wire [21:0] tlb_io_rent_ppn; // @[MMU.scala 65:19]
  wire  tlb_io_rent_d; // @[MMU.scala 65:19]
  wire  tlb_io_rent_a; // @[MMU.scala 65:19]
  wire  tlb_io_rent_u; // @[MMU.scala 65:19]
  wire  tlb_io_rent_x; // @[MMU.scala 65:19]
  wire  tlb_io_rent_w; // @[MMU.scala 65:19]
  wire  tlb_io_rent_r; // @[MMU.scala 65:19]
  reg [2:0] state; // @[MMU.scala 56:22]
  reg [31:0] _RAND_0;
  reg [21:0] entry_ppn; // @[MMU.scala 59:18]
  reg [31:0] _RAND_1;
  reg  entry_d; // @[MMU.scala 59:18]
  reg [31:0] _RAND_2;
  reg  entry_a; // @[MMU.scala 59:18]
  reg [31:0] _RAND_3;
  reg  entry_u; // @[MMU.scala 59:18]
  reg [31:0] _RAND_4;
  reg  entry_x; // @[MMU.scala 59:18]
  reg [31:0] _RAND_5;
  reg  entry_w; // @[MMU.scala 59:18]
  reg [31:0] _RAND_6;
  reg  entry_r; // @[MMU.scala 59:18]
  reg [31:0] _RAND_7;
  reg [31:0] addr; // @[MMU.scala 60:18]
  reg [31:0] _RAND_8;
  reg  level; // @[MMU.scala 61:18]
  reg [31:0] _RAND_9;
  wire  pte_v = io_data_rdata[0]; // @[MMU.scala 62:55]
  wire  pte_r = io_data_rdata[1]; // @[MMU.scala 62:55]
  wire  pte_w = io_data_rdata[2]; // @[MMU.scala 62:55]
  wire  pte_x = io_data_rdata[3]; // @[MMU.scala 62:55]
  wire  pte_u = io_data_rdata[4]; // @[MMU.scala 62:55]
  wire  pte_a = io_data_rdata[6]; // @[MMU.scala 62:55]
  wire  pte_d = io_data_rdata[7]; // @[MMU.scala 62:55]
  wire [21:0] pte_ppn = io_data_rdata[31:10]; // @[MMU.scala 62:55]
  wire  tlbFlush = state == 3'h4; // @[MMU.scala 72:25]
  wire  _T_13 = state == 3'h0; // @[MMU.scala 73:25]
  wire  tlbHit = _T_13 & tlb_io_valid; // @[MMU.scala 73:35]
  wire  _T_14 = ~io_en; // @[MMU.scala 74:19]
  wire  _T_15 = _T_14 | tlbFlush; // @[MMU.scala 74:26]
  wire  valid = _T_15 | tlbHit; // @[MMU.scala 74:38]
  wire  daFault = ~tlb_io_rent_a; // @[MMU.scala 77:17]
  wire  xFault = ~tlb_io_rent_x; // @[MMU.scala 80:29]
  wire  _T_20 = ~io_sum; // @[MMU.scala 81:29]
  wire  _T_21 = io_smode & _T_20; // @[MMU.scala 81:26]
  wire  uFault = _T_21 & tlb_io_rent_u; // @[MMU.scala 81:37]
  wire  _T_24 = daFault | xFault; // @[MMU.scala 82:45]
  wire  vmFault = _T_24 | uFault; // @[MMU.scala 82:55]
  wire  fault = io_en & vmFault; // @[MMU.scala 83:23]
  wire [11:0] voffset = io_vaddr[11:0]; // @[MMU.scala 86:25]
  wire [33:0] _T_25 = {tlb_io_rent_ppn,voffset}; // @[Cat.scala 30:58]
  wire [31:0] tlbAddr = _T_25[31:0]; // @[MMU.scala 87:46]
  wire  _T_26 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_27 = ~tlb_io_valid; // @[MMU.scala 103:28]
  wire [33:0] _T_29 = {io_basePpn, 12'h0}; // @[Paging.scala 41:12]
  wire [11:0] _T_34 = {io_vaddr[31:22], 2'h0}; // @[Paging.scala 41:51]
  wire [33:0] _GEN_82 = {{22'd0}, _T_34}; // @[Paging.scala 41:27]
  wire [33:0] _T_36 = _T_29 + _GEN_82; // @[Paging.scala 41:27]
  wire [33:0] _GEN_1 = _T_27 ? _T_36 : {{2'd0}, addr}; // @[MMU.scala 103:43]
  wire  _GEN_2 = _T_27 | level; // @[MMU.scala 103:43]
  wire [33:0] _GEN_4 = io_en ? _GEN_1 : {{2'd0}, addr}; // @[MMU.scala 101:27]
  wire [33:0] _GEN_7 = io_flush ? {{2'd0}, addr} : _GEN_4; // @[MMU.scala 98:23]
  wire  _T_37 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_38 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_39 = ~pte_v; // @[MMU.scala 118:13]
  wire  _T_40 = ~pte_r; // @[MMU.scala 118:24]
  wire  _T_41 = _T_40 & pte_w; // @[MMU.scala 118:31]
  wire  _T_42 = _T_39 | _T_41; // @[MMU.scala 118:20]
  wire  _T_44 = pte_r | pte_x; // @[MMU.scala 121:26]
  wire  _T_45 = level > 1'h0; // @[MMU.scala 122:21]
  wire  _T_47 = level - 1'h1; // @[MMU.scala 122:58]
  wire [21:0] _T_51 = _T_47 ? pte_ppn : {{12'd0}, pte_ppn[9:0]}; // @[Paging.scala 37:10]
  wire  _T_52 = _T_51 != 22'h0; // @[MMU.scala 122:65]
  wire  _T_53 = _T_45 & _T_52; // @[MMU.scala 122:27]
  wire [21:0] _T_63 = pte_ppn ^ _T_51; // @[Paging.scala 45:12]
  wire [19:0] _T_67 = _T_47 ? io_vaddr[31:12] : {{10'd0}, io_vaddr[21:12]}; // @[Paging.scala 29:10]
  wire [21:0] _GEN_83 = {{2'd0}, _T_67}; // @[Paging.scala 45:40]
  wire [21:0] _T_68 = _T_63 | _GEN_83; // @[Paging.scala 45:40]
  wire  _T_69 = ~level; // @[MMU.scala 134:26]
  wire [33:0] _T_73 = {pte_ppn, 12'h0}; // @[Paging.scala 41:12]
  wire [9:0] _T_77 = _T_47 ? io_vaddr[31:22] : io_vaddr[21:12]; // @[Paging.scala 25:10]
  wire [11:0] _T_78 = {_T_77, 2'h0}; // @[Paging.scala 41:51]
  wire [33:0] _GEN_84 = {{22'd0}, _T_78}; // @[Paging.scala 41:27]
  wire [33:0] _T_80 = _T_73 + _GEN_84; // @[Paging.scala 41:27]
  wire [33:0] _GEN_27 = _T_69 ? {{2'd0}, addr} : _T_80; // @[MMU.scala 134:35]
  wire [33:0] _GEN_37 = _T_44 ? {{2'd0}, addr} : _GEN_27; // @[MMU.scala 121:36]
  wire [33:0] _GEN_47 = _T_42 ? {{2'd0}, addr} : _GEN_37; // @[MMU.scala 118:42]
  wire  _T_83 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_84 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_85 = ~io_flush; // @[MMU.scala 150:13]
  wire [33:0] _GEN_60 = _T_38 ? _GEN_47 : {{2'd0}, addr}; // @[Conditional.scala 39:67]
  wire [33:0] _GEN_70 = _T_37 ? {{2'd0}, addr} : _GEN_60; // @[Conditional.scala 39:67]
  wire [33:0] _GEN_73 = _T_26 ? _GEN_7 : _GEN_70; // @[Conditional.scala 40:58]
  TLB tlb ( // @[MMU.scala 65:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_flush(tlb_io_flush),
    .io_wen(tlb_io_wen),
    .io_vaddr(tlb_io_vaddr),
    .io_went_ppn(tlb_io_went_ppn),
    .io_went_d(tlb_io_went_d),
    .io_went_a(tlb_io_went_a),
    .io_went_u(tlb_io_went_u),
    .io_went_x(tlb_io_went_x),
    .io_went_w(tlb_io_went_w),
    .io_went_r(tlb_io_went_r),
    .io_valid(tlb_io_valid),
    .io_rent_ppn(tlb_io_rent_ppn),
    .io_rent_d(tlb_io_rent_d),
    .io_rent_a(tlb_io_rent_a),
    .io_rent_u(tlb_io_rent_u),
    .io_rent_x(tlb_io_rent_x),
    .io_rent_w(tlb_io_rent_w),
    .io_rent_r(tlb_io_rent_r)
  );
  assign io_valid = _T_15 | tlbHit; // @[MMU.scala 161:13]
  assign io_fault = valid & fault; // @[MMU.scala 162:13]
  assign io_paddr = io_en ? tlbAddr : io_vaddr; // @[MMU.scala 163:13]
  assign io_data_en = state == 3'h1; // @[MMU.scala 155:17]
  assign io_data_addr = addr; // @[MMU.scala 157:17]
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_flush = io_flush; // @[MMU.scala 66:17]
  assign tlb_io_wen = state == 3'h3; // @[MMU.scala 67:17]
  assign tlb_io_vaddr = io_vaddr; // @[MMU.scala 68:17]
  assign tlb_io_went_ppn = entry_ppn; // @[MMU.scala 69:17]
  assign tlb_io_went_d = entry_d; // @[MMU.scala 69:17]
  assign tlb_io_went_a = entry_a; // @[MMU.scala 69:17]
  assign tlb_io_went_u = entry_u; // @[MMU.scala 69:17]
  assign tlb_io_went_x = entry_x; // @[MMU.scala 69:17]
  assign tlb_io_went_w = entry_w; // @[MMU.scala 69:17]
  assign tlb_io_went_r = entry_r; // @[MMU.scala 69:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  entry_ppn = _RAND_1[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  entry_d = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  entry_a = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  entry_u = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  entry_x = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  entry_w = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  entry_r = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  level = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (_T_26) begin
      if (io_flush) begin
        state <= 3'h4;
      end else if (io_en) begin
        if (_T_27) begin
          state <= 3'h1;
        end
      end
    end else if (_T_37) begin
      if (io_data_valid) begin
        state <= 3'h2;
      end
    end else if (_T_38) begin
      if (_T_42) begin
        state <= 3'h3;
      end else if (_T_44) begin
        state <= 3'h3;
      end else if (_T_69) begin
        state <= 3'h3;
      end else begin
        state <= 3'h1;
      end
    end else if (_T_83) begin
      state <= 3'h0;
    end else if (_T_84) begin
      if (_T_85) begin
        state <= 3'h0;
      end
    end
    if (!(_T_26)) begin
      if (!(_T_37)) begin
        if (_T_38) begin
          if (_T_42) begin
            entry_ppn <= 22'h0;
          end else if (_T_44) begin
            if (_T_53) begin
              entry_ppn <= 22'h0;
            end else if (_T_45) begin
              entry_ppn <= _T_68;
            end else begin
              entry_ppn <= pte_ppn;
            end
          end else if (_T_69) begin
            entry_ppn <= 22'h0;
          end
        end
      end
    end
    if (!(_T_26)) begin
      if (!(_T_37)) begin
        if (_T_38) begin
          if (_T_42) begin
            entry_d <= 1'h0;
          end else if (_T_44) begin
            if (_T_53) begin
              entry_d <= 1'h0;
            end else begin
              entry_d <= pte_d;
            end
          end else if (_T_69) begin
            entry_d <= 1'h0;
          end
        end
      end
    end
    if (!(_T_26)) begin
      if (!(_T_37)) begin
        if (_T_38) begin
          if (_T_42) begin
            entry_a <= 1'h0;
          end else if (_T_44) begin
            if (_T_53) begin
              entry_a <= 1'h0;
            end else begin
              entry_a <= pte_a;
            end
          end else if (_T_69) begin
            entry_a <= 1'h0;
          end
        end
      end
    end
    if (!(_T_26)) begin
      if (!(_T_37)) begin
        if (_T_38) begin
          if (_T_42) begin
            entry_u <= 1'h0;
          end else if (_T_44) begin
            if (_T_53) begin
              entry_u <= 1'h0;
            end else begin
              entry_u <= pte_u;
            end
          end else if (_T_69) begin
            entry_u <= 1'h0;
          end
        end
      end
    end
    if (!(_T_26)) begin
      if (!(_T_37)) begin
        if (_T_38) begin
          if (_T_42) begin
            entry_x <= 1'h0;
          end else if (_T_44) begin
            if (_T_53) begin
              entry_x <= 1'h0;
            end else begin
              entry_x <= pte_x;
            end
          end else if (_T_69) begin
            entry_x <= 1'h0;
          end
        end
      end
    end
    if (!(_T_26)) begin
      if (!(_T_37)) begin
        if (_T_38) begin
          if (_T_42) begin
            entry_w <= 1'h0;
          end else if (_T_44) begin
            if (_T_53) begin
              entry_w <= 1'h0;
            end else begin
              entry_w <= pte_w;
            end
          end else if (_T_69) begin
            entry_w <= 1'h0;
          end
        end
      end
    end
    if (!(_T_26)) begin
      if (!(_T_37)) begin
        if (_T_38) begin
          if (_T_42) begin
            entry_r <= 1'h0;
          end else if (_T_44) begin
            if (_T_53) begin
              entry_r <= 1'h0;
            end else begin
              entry_r <= pte_r;
            end
          end else if (_T_69) begin
            entry_r <= 1'h0;
          end
        end
      end
    end
    addr <= _GEN_73[31:0];
    if (_T_26) begin
      if (!(io_flush)) begin
        if (io_en) begin
          level <= _GEN_2;
        end
      end
    end else if (!(_T_37)) begin
      if (_T_38) begin
        if (!(_T_42)) begin
          if (!(_T_44)) begin
            if (!(_T_69)) begin
              level <= _T_47;
            end
          end
        end
      end
    end
  end
endmodule
module SramDemux2(
  input         io_sel2,
  input         io_in1_en,
  output        io_in1_valid,
  input  [31:0] io_in1_addr,
  output [31:0] io_in1_rdata,
  input         io_in2_en,
  output        io_in2_valid,
  input  [3:0]  io_in2_wen,
  input  [31:0] io_in2_addr,
  output [31:0] io_in2_rdata,
  input  [31:0] io_in2_wdata,
  output        io_out_en,
  input         io_out_valid,
  output [3:0]  io_out_wen,
  output [31:0] io_out_addr,
  input  [31:0] io_out_rdata,
  output [31:0] io_out_wdata
);
  wire  _T = ~io_sel2; // @[SramUtils.scala 41:20]
  assign io_in1_valid = _T & io_out_valid; // @[SramUtils.scala 41:17]
  assign io_in1_rdata = io_out_rdata; // @[SramUtils.scala 43:17]
  assign io_in2_valid = io_sel2 & io_out_valid; // @[SramUtils.scala 45:17]
  assign io_in2_rdata = io_out_rdata; // @[SramUtils.scala 47:17]
  assign io_out_en = io_sel2 ? io_in2_en : io_in1_en; // @[SramUtils.scala 49:17]
  assign io_out_wen = io_sel2 ? io_in2_wen : 4'h0; // @[SramUtils.scala 50:17]
  assign io_out_addr = io_sel2 ? io_in2_addr : io_in1_addr; // @[SramUtils.scala 51:17]
  assign io_out_wdata = io_sel2 ? io_in2_wdata : 32'h0; // @[SramUtils.scala 52:17]
endmodule
module InstCache(
  input         clock,
  input         reset,
  input         io_sram_en,
  output        io_sram_valid,
  input  [31:0] io_sram_addr,
  output [31:0] io_sram_rdata,
  input         io_flush,
  input         io_axi_readAddr_ready,
  output        io_axi_readAddr_valid,
  output [31:0] io_axi_readAddr_bits_addr,
  input         io_axi_readData_valid,
  input  [31:0] io_axi_readData_bits_data,
  input         io_axi_readData_bits_last
);
  reg [19:0] tag [0:63]; // @[InstCache.scala 34:18]
  reg [31:0] _RAND_0;
  wire [19:0] tag__T_3_data; // @[InstCache.scala 34:18]
  wire [5:0] tag__T_3_addr; // @[InstCache.scala 34:18]
  wire [19:0] tag__T_15_data; // @[InstCache.scala 34:18]
  wire [5:0] tag__T_15_addr; // @[InstCache.scala 34:18]
  wire  tag__T_15_mask; // @[InstCache.scala 34:18]
  wire  tag__T_15_en; // @[InstCache.scala 34:18]
  reg [31:0] lines [0:1023]; // @[InstCache.scala 35:26]
  reg [31:0] _RAND_1;
  wire [31:0] lines__T_18_data; // @[InstCache.scala 35:26]
  wire [9:0] lines__T_18_addr; // @[InstCache.scala 35:26]
  wire [31:0] lines__T_12_data; // @[InstCache.scala 35:26]
  wire [9:0] lines__T_12_addr; // @[InstCache.scala 35:26]
  wire  lines__T_12_mask; // @[InstCache.scala 35:26]
  wire  lines__T_12_en; // @[InstCache.scala 35:26]
  reg  lines__T_18_en_pipe_0;
  reg [31:0] _RAND_2;
  reg [9:0] lines__T_18_addr_pipe_0;
  reg [31:0] _RAND_3;
  reg [1:0] state; // @[InstCache.scala 30:22]
  reg [31:0] _RAND_4;
  reg  valid_0; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_5;
  reg  valid_1; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_6;
  reg  valid_2; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_7;
  reg  valid_3; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_8;
  reg  valid_4; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_9;
  reg  valid_5; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_10;
  reg  valid_6; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_11;
  reg  valid_7; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_12;
  reg  valid_8; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_13;
  reg  valid_9; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_14;
  reg  valid_10; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_15;
  reg  valid_11; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_16;
  reg  valid_12; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_17;
  reg  valid_13; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_18;
  reg  valid_14; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_19;
  reg  valid_15; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_20;
  reg  valid_16; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_21;
  reg  valid_17; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_22;
  reg  valid_18; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_23;
  reg  valid_19; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_24;
  reg  valid_20; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_25;
  reg  valid_21; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_26;
  reg  valid_22; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_27;
  reg  valid_23; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_28;
  reg  valid_24; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_29;
  reg  valid_25; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_30;
  reg  valid_26; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_31;
  reg  valid_27; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_32;
  reg  valid_28; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_33;
  reg  valid_29; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_34;
  reg  valid_30; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_35;
  reg  valid_31; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_36;
  reg  valid_32; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_37;
  reg  valid_33; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_38;
  reg  valid_34; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_39;
  reg  valid_35; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_40;
  reg  valid_36; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_41;
  reg  valid_37; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_42;
  reg  valid_38; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_43;
  reg  valid_39; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_44;
  reg  valid_40; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_45;
  reg  valid_41; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_46;
  reg  valid_42; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_47;
  reg  valid_43; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_48;
  reg  valid_44; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_49;
  reg  valid_45; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_50;
  reg  valid_46; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_51;
  reg  valid_47; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_52;
  reg  valid_48; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_53;
  reg  valid_49; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_54;
  reg  valid_50; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_55;
  reg  valid_51; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_56;
  reg  valid_52; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_57;
  reg  valid_53; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_58;
  reg  valid_54; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_59;
  reg  valid_55; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_60;
  reg  valid_56; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_61;
  reg  valid_57; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_62;
  reg  valid_58; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_63;
  reg  valid_59; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_64;
  reg  valid_60; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_65;
  reg  valid_61; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_66;
  reg  valid_62; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_67;
  reg  valid_63; // @[InstCache.scala 33:22]
  reg [31:0] _RAND_68;
  reg  ren; // @[InstCache.scala 38:28]
  reg [31:0] _RAND_69;
  reg [31:0] raddr; // @[InstCache.scala 39:24]
  reg [31:0] _RAND_70;
  reg [3:0] dataOffset; // @[InstCache.scala 40:24]
  reg [31:0] _RAND_71;
  reg [31:0] sramAddr; // @[InstCache.scala 43:24]
  reg [31:0] _RAND_72;
  wire  _T_1 = state == 2'h0; // @[InstCache.scala 44:31]
  wire [31:0] selAddr = _T_1 ? io_sram_addr : sramAddr; // @[InstCache.scala 44:24]
  wire [19:0] tagSel = selAddr[31:12]; // @[InstCache.scala 45:28]
  wire [5:0] lineSel = selAddr[11:6]; // @[InstCache.scala 47:28]
  wire [31:0] startAddr = {tagSel,lineSel,6'h0}; // @[Cat.scala 30:58]
  wire  _T_4 = tag__T_3_data == tagSel; // @[InstCache.scala 53:52]
  wire  _GEN_1 = 6'h1 == lineSel ? valid_1 : valid_0; // @[InstCache.scala 53:36]
  wire  _GEN_2 = 6'h2 == lineSel ? valid_2 : _GEN_1; // @[InstCache.scala 53:36]
  wire  _GEN_3 = 6'h3 == lineSel ? valid_3 : _GEN_2; // @[InstCache.scala 53:36]
  wire  _GEN_4 = 6'h4 == lineSel ? valid_4 : _GEN_3; // @[InstCache.scala 53:36]
  wire  _GEN_5 = 6'h5 == lineSel ? valid_5 : _GEN_4; // @[InstCache.scala 53:36]
  wire  _GEN_6 = 6'h6 == lineSel ? valid_6 : _GEN_5; // @[InstCache.scala 53:36]
  wire  _GEN_7 = 6'h7 == lineSel ? valid_7 : _GEN_6; // @[InstCache.scala 53:36]
  wire  _GEN_8 = 6'h8 == lineSel ? valid_8 : _GEN_7; // @[InstCache.scala 53:36]
  wire  _GEN_9 = 6'h9 == lineSel ? valid_9 : _GEN_8; // @[InstCache.scala 53:36]
  wire  _GEN_10 = 6'ha == lineSel ? valid_10 : _GEN_9; // @[InstCache.scala 53:36]
  wire  _GEN_11 = 6'hb == lineSel ? valid_11 : _GEN_10; // @[InstCache.scala 53:36]
  wire  _GEN_12 = 6'hc == lineSel ? valid_12 : _GEN_11; // @[InstCache.scala 53:36]
  wire  _GEN_13 = 6'hd == lineSel ? valid_13 : _GEN_12; // @[InstCache.scala 53:36]
  wire  _GEN_14 = 6'he == lineSel ? valid_14 : _GEN_13; // @[InstCache.scala 53:36]
  wire  _GEN_15 = 6'hf == lineSel ? valid_15 : _GEN_14; // @[InstCache.scala 53:36]
  wire  _GEN_16 = 6'h10 == lineSel ? valid_16 : _GEN_15; // @[InstCache.scala 53:36]
  wire  _GEN_17 = 6'h11 == lineSel ? valid_17 : _GEN_16; // @[InstCache.scala 53:36]
  wire  _GEN_18 = 6'h12 == lineSel ? valid_18 : _GEN_17; // @[InstCache.scala 53:36]
  wire  _GEN_19 = 6'h13 == lineSel ? valid_19 : _GEN_18; // @[InstCache.scala 53:36]
  wire  _GEN_20 = 6'h14 == lineSel ? valid_20 : _GEN_19; // @[InstCache.scala 53:36]
  wire  _GEN_21 = 6'h15 == lineSel ? valid_21 : _GEN_20; // @[InstCache.scala 53:36]
  wire  _GEN_22 = 6'h16 == lineSel ? valid_22 : _GEN_21; // @[InstCache.scala 53:36]
  wire  _GEN_23 = 6'h17 == lineSel ? valid_23 : _GEN_22; // @[InstCache.scala 53:36]
  wire  _GEN_24 = 6'h18 == lineSel ? valid_24 : _GEN_23; // @[InstCache.scala 53:36]
  wire  _GEN_25 = 6'h19 == lineSel ? valid_25 : _GEN_24; // @[InstCache.scala 53:36]
  wire  _GEN_26 = 6'h1a == lineSel ? valid_26 : _GEN_25; // @[InstCache.scala 53:36]
  wire  _GEN_27 = 6'h1b == lineSel ? valid_27 : _GEN_26; // @[InstCache.scala 53:36]
  wire  _GEN_28 = 6'h1c == lineSel ? valid_28 : _GEN_27; // @[InstCache.scala 53:36]
  wire  _GEN_29 = 6'h1d == lineSel ? valid_29 : _GEN_28; // @[InstCache.scala 53:36]
  wire  _GEN_30 = 6'h1e == lineSel ? valid_30 : _GEN_29; // @[InstCache.scala 53:36]
  wire  _GEN_31 = 6'h1f == lineSel ? valid_31 : _GEN_30; // @[InstCache.scala 53:36]
  wire  _GEN_32 = 6'h20 == lineSel ? valid_32 : _GEN_31; // @[InstCache.scala 53:36]
  wire  _GEN_33 = 6'h21 == lineSel ? valid_33 : _GEN_32; // @[InstCache.scala 53:36]
  wire  _GEN_34 = 6'h22 == lineSel ? valid_34 : _GEN_33; // @[InstCache.scala 53:36]
  wire  _GEN_35 = 6'h23 == lineSel ? valid_35 : _GEN_34; // @[InstCache.scala 53:36]
  wire  _GEN_36 = 6'h24 == lineSel ? valid_36 : _GEN_35; // @[InstCache.scala 53:36]
  wire  _GEN_37 = 6'h25 == lineSel ? valid_37 : _GEN_36; // @[InstCache.scala 53:36]
  wire  _GEN_38 = 6'h26 == lineSel ? valid_38 : _GEN_37; // @[InstCache.scala 53:36]
  wire  _GEN_39 = 6'h27 == lineSel ? valid_39 : _GEN_38; // @[InstCache.scala 53:36]
  wire  _GEN_40 = 6'h28 == lineSel ? valid_40 : _GEN_39; // @[InstCache.scala 53:36]
  wire  _GEN_41 = 6'h29 == lineSel ? valid_41 : _GEN_40; // @[InstCache.scala 53:36]
  wire  _GEN_42 = 6'h2a == lineSel ? valid_42 : _GEN_41; // @[InstCache.scala 53:36]
  wire  _GEN_43 = 6'h2b == lineSel ? valid_43 : _GEN_42; // @[InstCache.scala 53:36]
  wire  _GEN_44 = 6'h2c == lineSel ? valid_44 : _GEN_43; // @[InstCache.scala 53:36]
  wire  _GEN_45 = 6'h2d == lineSel ? valid_45 : _GEN_44; // @[InstCache.scala 53:36]
  wire  _GEN_46 = 6'h2e == lineSel ? valid_46 : _GEN_45; // @[InstCache.scala 53:36]
  wire  _GEN_47 = 6'h2f == lineSel ? valid_47 : _GEN_46; // @[InstCache.scala 53:36]
  wire  _GEN_48 = 6'h30 == lineSel ? valid_48 : _GEN_47; // @[InstCache.scala 53:36]
  wire  _GEN_49 = 6'h31 == lineSel ? valid_49 : _GEN_48; // @[InstCache.scala 53:36]
  wire  _GEN_50 = 6'h32 == lineSel ? valid_50 : _GEN_49; // @[InstCache.scala 53:36]
  wire  _GEN_51 = 6'h33 == lineSel ? valid_51 : _GEN_50; // @[InstCache.scala 53:36]
  wire  _GEN_52 = 6'h34 == lineSel ? valid_52 : _GEN_51; // @[InstCache.scala 53:36]
  wire  _GEN_53 = 6'h35 == lineSel ? valid_53 : _GEN_52; // @[InstCache.scala 53:36]
  wire  _GEN_54 = 6'h36 == lineSel ? valid_54 : _GEN_53; // @[InstCache.scala 53:36]
  wire  _GEN_55 = 6'h37 == lineSel ? valid_55 : _GEN_54; // @[InstCache.scala 53:36]
  wire  _GEN_56 = 6'h38 == lineSel ? valid_56 : _GEN_55; // @[InstCache.scala 53:36]
  wire  _GEN_57 = 6'h39 == lineSel ? valid_57 : _GEN_56; // @[InstCache.scala 53:36]
  wire  _GEN_58 = 6'h3a == lineSel ? valid_58 : _GEN_57; // @[InstCache.scala 53:36]
  wire  _GEN_59 = 6'h3b == lineSel ? valid_59 : _GEN_58; // @[InstCache.scala 53:36]
  wire  _GEN_60 = 6'h3c == lineSel ? valid_60 : _GEN_59; // @[InstCache.scala 53:36]
  wire  _GEN_61 = 6'h3d == lineSel ? valid_61 : _GEN_60; // @[InstCache.scala 53:36]
  wire  _GEN_62 = 6'h3e == lineSel ? valid_62 : _GEN_61; // @[InstCache.scala 53:36]
  wire  _GEN_63 = 6'h3f == lineSel ? valid_63 : _GEN_62; // @[InstCache.scala 53:36]
  wire  cacheHit = _GEN_63 & _T_4; // @[InstCache.scala 53:36]
  wire  _T_5 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = ~cacheHit; // @[InstCache.scala 64:34]
  wire  _T_7 = io_sram_en & _T_6; // @[InstCache.scala 64:31]
  wire  _GEN_64 = _T_7 | ren; // @[InstCache.scala 64:45]
  wire  _T_8 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_9 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire [3:0] _T_11 = dataOffset + 4'h1; // @[InstCache.scala 84:34]
  wire  _T_13 = io_axi_readData_valid & io_axi_readData_bits_last; // @[InstCache.scala 88:35]
  wire  _T_14 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire  _GEN_512 = 6'h0 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_146 = _GEN_512 | valid_0; // @[InstCache.scala 94:23]
  wire  _GEN_513 = 6'h1 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_147 = _GEN_513 | valid_1; // @[InstCache.scala 94:23]
  wire  _GEN_514 = 6'h2 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_148 = _GEN_514 | valid_2; // @[InstCache.scala 94:23]
  wire  _GEN_515 = 6'h3 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_149 = _GEN_515 | valid_3; // @[InstCache.scala 94:23]
  wire  _GEN_516 = 6'h4 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_150 = _GEN_516 | valid_4; // @[InstCache.scala 94:23]
  wire  _GEN_517 = 6'h5 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_151 = _GEN_517 | valid_5; // @[InstCache.scala 94:23]
  wire  _GEN_518 = 6'h6 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_152 = _GEN_518 | valid_6; // @[InstCache.scala 94:23]
  wire  _GEN_519 = 6'h7 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_153 = _GEN_519 | valid_7; // @[InstCache.scala 94:23]
  wire  _GEN_520 = 6'h8 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_154 = _GEN_520 | valid_8; // @[InstCache.scala 94:23]
  wire  _GEN_521 = 6'h9 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_155 = _GEN_521 | valid_9; // @[InstCache.scala 94:23]
  wire  _GEN_522 = 6'ha == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_156 = _GEN_522 | valid_10; // @[InstCache.scala 94:23]
  wire  _GEN_523 = 6'hb == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_157 = _GEN_523 | valid_11; // @[InstCache.scala 94:23]
  wire  _GEN_524 = 6'hc == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_158 = _GEN_524 | valid_12; // @[InstCache.scala 94:23]
  wire  _GEN_525 = 6'hd == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_159 = _GEN_525 | valid_13; // @[InstCache.scala 94:23]
  wire  _GEN_526 = 6'he == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_160 = _GEN_526 | valid_14; // @[InstCache.scala 94:23]
  wire  _GEN_527 = 6'hf == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_161 = _GEN_527 | valid_15; // @[InstCache.scala 94:23]
  wire  _GEN_528 = 6'h10 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_162 = _GEN_528 | valid_16; // @[InstCache.scala 94:23]
  wire  _GEN_529 = 6'h11 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_163 = _GEN_529 | valid_17; // @[InstCache.scala 94:23]
  wire  _GEN_530 = 6'h12 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_164 = _GEN_530 | valid_18; // @[InstCache.scala 94:23]
  wire  _GEN_531 = 6'h13 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_165 = _GEN_531 | valid_19; // @[InstCache.scala 94:23]
  wire  _GEN_532 = 6'h14 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_166 = _GEN_532 | valid_20; // @[InstCache.scala 94:23]
  wire  _GEN_533 = 6'h15 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_167 = _GEN_533 | valid_21; // @[InstCache.scala 94:23]
  wire  _GEN_534 = 6'h16 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_168 = _GEN_534 | valid_22; // @[InstCache.scala 94:23]
  wire  _GEN_535 = 6'h17 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_169 = _GEN_535 | valid_23; // @[InstCache.scala 94:23]
  wire  _GEN_536 = 6'h18 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_170 = _GEN_536 | valid_24; // @[InstCache.scala 94:23]
  wire  _GEN_537 = 6'h19 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_171 = _GEN_537 | valid_25; // @[InstCache.scala 94:23]
  wire  _GEN_538 = 6'h1a == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_172 = _GEN_538 | valid_26; // @[InstCache.scala 94:23]
  wire  _GEN_539 = 6'h1b == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_173 = _GEN_539 | valid_27; // @[InstCache.scala 94:23]
  wire  _GEN_540 = 6'h1c == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_174 = _GEN_540 | valid_28; // @[InstCache.scala 94:23]
  wire  _GEN_541 = 6'h1d == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_175 = _GEN_541 | valid_29; // @[InstCache.scala 94:23]
  wire  _GEN_542 = 6'h1e == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_176 = _GEN_542 | valid_30; // @[InstCache.scala 94:23]
  wire  _GEN_543 = 6'h1f == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_177 = _GEN_543 | valid_31; // @[InstCache.scala 94:23]
  wire  _GEN_544 = 6'h20 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_178 = _GEN_544 | valid_32; // @[InstCache.scala 94:23]
  wire  _GEN_545 = 6'h21 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_179 = _GEN_545 | valid_33; // @[InstCache.scala 94:23]
  wire  _GEN_546 = 6'h22 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_180 = _GEN_546 | valid_34; // @[InstCache.scala 94:23]
  wire  _GEN_547 = 6'h23 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_181 = _GEN_547 | valid_35; // @[InstCache.scala 94:23]
  wire  _GEN_548 = 6'h24 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_182 = _GEN_548 | valid_36; // @[InstCache.scala 94:23]
  wire  _GEN_549 = 6'h25 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_183 = _GEN_549 | valid_37; // @[InstCache.scala 94:23]
  wire  _GEN_550 = 6'h26 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_184 = _GEN_550 | valid_38; // @[InstCache.scala 94:23]
  wire  _GEN_551 = 6'h27 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_185 = _GEN_551 | valid_39; // @[InstCache.scala 94:23]
  wire  _GEN_552 = 6'h28 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_186 = _GEN_552 | valid_40; // @[InstCache.scala 94:23]
  wire  _GEN_553 = 6'h29 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_187 = _GEN_553 | valid_41; // @[InstCache.scala 94:23]
  wire  _GEN_554 = 6'h2a == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_188 = _GEN_554 | valid_42; // @[InstCache.scala 94:23]
  wire  _GEN_555 = 6'h2b == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_189 = _GEN_555 | valid_43; // @[InstCache.scala 94:23]
  wire  _GEN_556 = 6'h2c == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_190 = _GEN_556 | valid_44; // @[InstCache.scala 94:23]
  wire  _GEN_557 = 6'h2d == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_191 = _GEN_557 | valid_45; // @[InstCache.scala 94:23]
  wire  _GEN_558 = 6'h2e == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_192 = _GEN_558 | valid_46; // @[InstCache.scala 94:23]
  wire  _GEN_559 = 6'h2f == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_193 = _GEN_559 | valid_47; // @[InstCache.scala 94:23]
  wire  _GEN_560 = 6'h30 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_194 = _GEN_560 | valid_48; // @[InstCache.scala 94:23]
  wire  _GEN_561 = 6'h31 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_195 = _GEN_561 | valid_49; // @[InstCache.scala 94:23]
  wire  _GEN_562 = 6'h32 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_196 = _GEN_562 | valid_50; // @[InstCache.scala 94:23]
  wire  _GEN_563 = 6'h33 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_197 = _GEN_563 | valid_51; // @[InstCache.scala 94:23]
  wire  _GEN_564 = 6'h34 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_198 = _GEN_564 | valid_52; // @[InstCache.scala 94:23]
  wire  _GEN_565 = 6'h35 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_199 = _GEN_565 | valid_53; // @[InstCache.scala 94:23]
  wire  _GEN_566 = 6'h36 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_200 = _GEN_566 | valid_54; // @[InstCache.scala 94:23]
  wire  _GEN_567 = 6'h37 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_201 = _GEN_567 | valid_55; // @[InstCache.scala 94:23]
  wire  _GEN_568 = 6'h38 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_202 = _GEN_568 | valid_56; // @[InstCache.scala 94:23]
  wire  _GEN_569 = 6'h39 == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_203 = _GEN_569 | valid_57; // @[InstCache.scala 94:23]
  wire  _GEN_570 = 6'h3a == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_204 = _GEN_570 | valid_58; // @[InstCache.scala 94:23]
  wire  _GEN_571 = 6'h3b == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_205 = _GEN_571 | valid_59; // @[InstCache.scala 94:23]
  wire  _GEN_572 = 6'h3c == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_206 = _GEN_572 | valid_60; // @[InstCache.scala 94:23]
  wire  _GEN_573 = 6'h3d == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_207 = _GEN_573 | valid_61; // @[InstCache.scala 94:23]
  wire  _GEN_574 = 6'h3e == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_208 = _GEN_574 | valid_62; // @[InstCache.scala 94:23]
  wire  _GEN_575 = 6'h3f == lineSel; // @[InstCache.scala 94:23]
  wire  _GEN_209 = _GEN_575 | valid_63; // @[InstCache.scala 94:23]
  wire  _GEN_283 = _T_9 & io_axi_readData_valid; // @[Conditional.scala 39:67]
  wire  _GEN_353 = _T_9 ? 1'h0 : _T_14; // @[Conditional.scala 39:67]
  wire  _GEN_361 = _T_8 ? 1'h0 : _GEN_283; // @[Conditional.scala 39:67]
  wire  _GEN_430 = _T_8 ? 1'h0 : _GEN_353; // @[Conditional.scala 39:67]
  assign tag__T_3_addr = selAddr[11:6];
  assign tag__T_3_data = tag[tag__T_3_addr]; // @[InstCache.scala 34:18]
  assign tag__T_15_data = selAddr[31:12];
  assign tag__T_15_addr = selAddr[11:6];
  assign tag__T_15_mask = 1'h1;
  assign tag__T_15_en = _T_5 ? 1'h0 : _GEN_430;
  assign lines__T_18_addr = lines__T_18_addr_pipe_0;
  assign lines__T_18_data = lines[lines__T_18_addr]; // @[InstCache.scala 35:26]
  assign lines__T_12_data = io_axi_readData_bits_data;
  assign lines__T_12_addr = {lineSel,dataOffset};
  assign lines__T_12_mask = 1'h1;
  assign lines__T_12_en = _T_5 ? 1'h0 : _GEN_361;
  assign io_sram_valid = _T_1 & cacheHit; // @[InstCache.scala 101:17]
  assign io_sram_rdata = lines__T_18_data; // @[InstCache.scala 103:17]
  assign io_axi_readAddr_valid = ren; // @[AXI.scala 56:20 InstCache.scala 107:31]
  assign io_axi_readAddr_bits_addr = raddr; // @[AXI.scala 9:21 InstCache.scala 108:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag[initvar] = _RAND_0[19:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    lines[initvar] = _RAND_1[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  lines__T_18_en_pipe_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  lines__T_18_addr_pipe_0 = _RAND_3[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  state = _RAND_4[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  valid_0 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  valid_1 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  valid_2 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  valid_3 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  valid_4 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  valid_5 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  valid_6 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  valid_7 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  valid_8 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  valid_9 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  valid_10 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  valid_11 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  valid_12 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  valid_13 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  valid_14 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valid_15 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  valid_16 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  valid_17 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  valid_18 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  valid_19 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  valid_20 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  valid_21 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  valid_22 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  valid_23 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  valid_24 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  valid_25 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  valid_26 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  valid_27 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  valid_28 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  valid_29 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  valid_30 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  valid_31 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  valid_32 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  valid_33 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  valid_34 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  valid_35 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  valid_36 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  valid_37 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  valid_38 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  valid_39 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  valid_40 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  valid_41 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  valid_42 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  valid_43 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  valid_44 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  valid_45 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  valid_46 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  valid_47 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  valid_48 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  valid_49 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  valid_50 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  valid_51 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  valid_52 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  valid_53 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  valid_54 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  valid_55 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  valid_56 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  valid_57 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  valid_58 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  valid_59 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  valid_60 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  valid_61 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  valid_62 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  valid_63 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  ren = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  raddr = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  dataOffset = _RAND_71[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  sramAddr = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tag__T_15_en & tag__T_15_mask) begin
      tag[tag__T_15_addr] <= tag__T_15_data; // @[InstCache.scala 34:18]
    end
    if(lines__T_12_en & lines__T_12_mask) begin
      lines[lines__T_12_addr] <= lines__T_12_data; // @[InstCache.scala 35:26]
    end
    lines__T_18_en_pipe_0 <= 1'h1;
    lines__T_18_addr_pipe_0 <= selAddr[11:2];
    if (reset) begin
      state <= 2'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        state <= 2'h0;
      end else if (_T_7) begin
        state <= 2'h1;
      end
    end else if (_T_8) begin
      if (io_axi_readAddr_ready) begin
        state <= 2'h2;
      end
    end else if (_T_9) begin
      if (_T_13) begin
        state <= 2'h3;
      end
    end else if (_T_14) begin
      state <= 2'h0;
    end
    if (reset) begin
      valid_0 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_0 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_0 <= _GEN_146;
        end
      end
    end
    if (reset) begin
      valid_1 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_1 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_1 <= _GEN_147;
        end
      end
    end
    if (reset) begin
      valid_2 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_2 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_2 <= _GEN_148;
        end
      end
    end
    if (reset) begin
      valid_3 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_3 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_3 <= _GEN_149;
        end
      end
    end
    if (reset) begin
      valid_4 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_4 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_4 <= _GEN_150;
        end
      end
    end
    if (reset) begin
      valid_5 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_5 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_5 <= _GEN_151;
        end
      end
    end
    if (reset) begin
      valid_6 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_6 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_6 <= _GEN_152;
        end
      end
    end
    if (reset) begin
      valid_7 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_7 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_7 <= _GEN_153;
        end
      end
    end
    if (reset) begin
      valid_8 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_8 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_8 <= _GEN_154;
        end
      end
    end
    if (reset) begin
      valid_9 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_9 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_9 <= _GEN_155;
        end
      end
    end
    if (reset) begin
      valid_10 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_10 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_10 <= _GEN_156;
        end
      end
    end
    if (reset) begin
      valid_11 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_11 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_11 <= _GEN_157;
        end
      end
    end
    if (reset) begin
      valid_12 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_12 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_12 <= _GEN_158;
        end
      end
    end
    if (reset) begin
      valid_13 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_13 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_13 <= _GEN_159;
        end
      end
    end
    if (reset) begin
      valid_14 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_14 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_14 <= _GEN_160;
        end
      end
    end
    if (reset) begin
      valid_15 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_15 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_15 <= _GEN_161;
        end
      end
    end
    if (reset) begin
      valid_16 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_16 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_16 <= _GEN_162;
        end
      end
    end
    if (reset) begin
      valid_17 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_17 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_17 <= _GEN_163;
        end
      end
    end
    if (reset) begin
      valid_18 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_18 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_18 <= _GEN_164;
        end
      end
    end
    if (reset) begin
      valid_19 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_19 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_19 <= _GEN_165;
        end
      end
    end
    if (reset) begin
      valid_20 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_20 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_20 <= _GEN_166;
        end
      end
    end
    if (reset) begin
      valid_21 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_21 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_21 <= _GEN_167;
        end
      end
    end
    if (reset) begin
      valid_22 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_22 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_22 <= _GEN_168;
        end
      end
    end
    if (reset) begin
      valid_23 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_23 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_23 <= _GEN_169;
        end
      end
    end
    if (reset) begin
      valid_24 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_24 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_24 <= _GEN_170;
        end
      end
    end
    if (reset) begin
      valid_25 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_25 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_25 <= _GEN_171;
        end
      end
    end
    if (reset) begin
      valid_26 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_26 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_26 <= _GEN_172;
        end
      end
    end
    if (reset) begin
      valid_27 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_27 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_27 <= _GEN_173;
        end
      end
    end
    if (reset) begin
      valid_28 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_28 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_28 <= _GEN_174;
        end
      end
    end
    if (reset) begin
      valid_29 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_29 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_29 <= _GEN_175;
        end
      end
    end
    if (reset) begin
      valid_30 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_30 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_30 <= _GEN_176;
        end
      end
    end
    if (reset) begin
      valid_31 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_31 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_31 <= _GEN_177;
        end
      end
    end
    if (reset) begin
      valid_32 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_32 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_32 <= _GEN_178;
        end
      end
    end
    if (reset) begin
      valid_33 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_33 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_33 <= _GEN_179;
        end
      end
    end
    if (reset) begin
      valid_34 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_34 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_34 <= _GEN_180;
        end
      end
    end
    if (reset) begin
      valid_35 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_35 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_35 <= _GEN_181;
        end
      end
    end
    if (reset) begin
      valid_36 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_36 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_36 <= _GEN_182;
        end
      end
    end
    if (reset) begin
      valid_37 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_37 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_37 <= _GEN_183;
        end
      end
    end
    if (reset) begin
      valid_38 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_38 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_38 <= _GEN_184;
        end
      end
    end
    if (reset) begin
      valid_39 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_39 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_39 <= _GEN_185;
        end
      end
    end
    if (reset) begin
      valid_40 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_40 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_40 <= _GEN_186;
        end
      end
    end
    if (reset) begin
      valid_41 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_41 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_41 <= _GEN_187;
        end
      end
    end
    if (reset) begin
      valid_42 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_42 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_42 <= _GEN_188;
        end
      end
    end
    if (reset) begin
      valid_43 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_43 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_43 <= _GEN_189;
        end
      end
    end
    if (reset) begin
      valid_44 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_44 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_44 <= _GEN_190;
        end
      end
    end
    if (reset) begin
      valid_45 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_45 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_45 <= _GEN_191;
        end
      end
    end
    if (reset) begin
      valid_46 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_46 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_46 <= _GEN_192;
        end
      end
    end
    if (reset) begin
      valid_47 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_47 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_47 <= _GEN_193;
        end
      end
    end
    if (reset) begin
      valid_48 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_48 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_48 <= _GEN_194;
        end
      end
    end
    if (reset) begin
      valid_49 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_49 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_49 <= _GEN_195;
        end
      end
    end
    if (reset) begin
      valid_50 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_50 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_50 <= _GEN_196;
        end
      end
    end
    if (reset) begin
      valid_51 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_51 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_51 <= _GEN_197;
        end
      end
    end
    if (reset) begin
      valid_52 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_52 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_52 <= _GEN_198;
        end
      end
    end
    if (reset) begin
      valid_53 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_53 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_53 <= _GEN_199;
        end
      end
    end
    if (reset) begin
      valid_54 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_54 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_54 <= _GEN_200;
        end
      end
    end
    if (reset) begin
      valid_55 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_55 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_55 <= _GEN_201;
        end
      end
    end
    if (reset) begin
      valid_56 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_56 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_56 <= _GEN_202;
        end
      end
    end
    if (reset) begin
      valid_57 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_57 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_57 <= _GEN_203;
        end
      end
    end
    if (reset) begin
      valid_58 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_58 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_58 <= _GEN_204;
        end
      end
    end
    if (reset) begin
      valid_59 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_59 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_59 <= _GEN_205;
        end
      end
    end
    if (reset) begin
      valid_60 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_60 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_60 <= _GEN_206;
        end
      end
    end
    if (reset) begin
      valid_61 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_61 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_61 <= _GEN_207;
        end
      end
    end
    if (reset) begin
      valid_62 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_62 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_62 <= _GEN_208;
        end
      end
    end
    if (reset) begin
      valid_63 <= 1'h0;
    end else if (_T_5) begin
      if (io_flush) begin
        valid_63 <= 1'h0;
      end
    end else if (!(_T_8)) begin
      if (!(_T_9)) begin
        if (_T_14) begin
          valid_63 <= _GEN_209;
        end
      end
    end
    if (reset) begin
      ren <= 1'h0;
    end else if (_T_5) begin
      if (!(io_flush)) begin
        ren <= _GEN_64;
      end
    end else if (_T_8) begin
      if (io_axi_readAddr_ready) begin
        ren <= 1'h0;
      end
    end
    if (_T_5) begin
      if (!(io_flush)) begin
        if (_T_7) begin
          raddr <= startAddr;
        end
      end
    end
    if (!(_T_5)) begin
      if (_T_8) begin
        if (io_axi_readAddr_ready) begin
          dataOffset <= 4'h0;
        end
      end else if (_T_9) begin
        if (io_axi_readData_valid) begin
          dataOffset <= _T_11;
        end
      end
    end
    if (_T_5) begin
      if (!(io_flush)) begin
        if (_T_7) begin
          sramAddr <= io_sram_addr;
        end
      end
    end
  end
endmodule
module MMU_1(
  input         clock,
  input         reset,
  input         io_en,
  input         io_flush,
  input  [21:0] io_basePpn,
  input         io_sum,
  input         io_smode,
  input         io_lookup,
  input         io_write,
  input  [31:0] io_vaddr,
  output        io_valid,
  output        io_fault,
  output [31:0] io_paddr,
  output        io_data_en,
  input         io_data_valid,
  output [31:0] io_data_addr,
  input  [31:0] io_data_rdata
);
  wire  tlb_clock; // @[MMU.scala 65:19]
  wire  tlb_reset; // @[MMU.scala 65:19]
  wire  tlb_io_flush; // @[MMU.scala 65:19]
  wire  tlb_io_wen; // @[MMU.scala 65:19]
  wire [31:0] tlb_io_vaddr; // @[MMU.scala 65:19]
  wire [21:0] tlb_io_went_ppn; // @[MMU.scala 65:19]
  wire  tlb_io_went_d; // @[MMU.scala 65:19]
  wire  tlb_io_went_a; // @[MMU.scala 65:19]
  wire  tlb_io_went_u; // @[MMU.scala 65:19]
  wire  tlb_io_went_x; // @[MMU.scala 65:19]
  wire  tlb_io_went_w; // @[MMU.scala 65:19]
  wire  tlb_io_went_r; // @[MMU.scala 65:19]
  wire  tlb_io_valid; // @[MMU.scala 65:19]
  wire [21:0] tlb_io_rent_ppn; // @[MMU.scala 65:19]
  wire  tlb_io_rent_d; // @[MMU.scala 65:19]
  wire  tlb_io_rent_a; // @[MMU.scala 65:19]
  wire  tlb_io_rent_u; // @[MMU.scala 65:19]
  wire  tlb_io_rent_x; // @[MMU.scala 65:19]
  wire  tlb_io_rent_w; // @[MMU.scala 65:19]
  wire  tlb_io_rent_r; // @[MMU.scala 65:19]
  reg [2:0] state; // @[MMU.scala 56:22]
  reg [31:0] _RAND_0;
  reg [21:0] entry_ppn; // @[MMU.scala 59:18]
  reg [31:0] _RAND_1;
  reg  entry_d; // @[MMU.scala 59:18]
  reg [31:0] _RAND_2;
  reg  entry_a; // @[MMU.scala 59:18]
  reg [31:0] _RAND_3;
  reg  entry_u; // @[MMU.scala 59:18]
  reg [31:0] _RAND_4;
  reg  entry_x; // @[MMU.scala 59:18]
  reg [31:0] _RAND_5;
  reg  entry_w; // @[MMU.scala 59:18]
  reg [31:0] _RAND_6;
  reg  entry_r; // @[MMU.scala 59:18]
  reg [31:0] _RAND_7;
  reg [31:0] addr; // @[MMU.scala 60:18]
  reg [31:0] _RAND_8;
  reg  level; // @[MMU.scala 61:18]
  reg [31:0] _RAND_9;
  wire  pte_v = io_data_rdata[0]; // @[MMU.scala 62:55]
  wire  pte_r = io_data_rdata[1]; // @[MMU.scala 62:55]
  wire  pte_w = io_data_rdata[2]; // @[MMU.scala 62:55]
  wire  pte_x = io_data_rdata[3]; // @[MMU.scala 62:55]
  wire  pte_u = io_data_rdata[4]; // @[MMU.scala 62:55]
  wire  pte_a = io_data_rdata[6]; // @[MMU.scala 62:55]
  wire  pte_d = io_data_rdata[7]; // @[MMU.scala 62:55]
  wire [21:0] pte_ppn = io_data_rdata[31:10]; // @[MMU.scala 62:55]
  wire  tlbFlush = state == 3'h4; // @[MMU.scala 72:25]
  wire  _T_13 = state == 3'h0; // @[MMU.scala 73:25]
  wire  tlbHit = _T_13 & tlb_io_valid; // @[MMU.scala 73:35]
  wire  _T_14 = ~io_en; // @[MMU.scala 74:19]
  wire  _T_15 = _T_14 | tlbFlush; // @[MMU.scala 74:26]
  wire  valid = _T_15 | tlbHit; // @[MMU.scala 74:38]
  wire  _T_16 = ~tlb_io_rent_a; // @[MMU.scala 77:17]
  wire  _T_17 = ~tlb_io_rent_d; // @[MMU.scala 77:48]
  wire  _T_18 = io_write & _T_17; // @[MMU.scala 77:45]
  wire  daFault = _T_16 | _T_18; // @[MMU.scala 77:32]
  wire  _T_19 = ~io_write; // @[MMU.scala 78:30]
  wire  _T_20 = ~tlb_io_rent_r; // @[MMU.scala 78:43]
  wire  rFault = _T_19 & _T_20; // @[MMU.scala 78:40]
  wire  _T_21 = ~tlb_io_rent_w; // @[MMU.scala 79:29]
  wire  wFault = io_write & _T_21; // @[MMU.scala 79:26]
  wire  _T_22 = ~io_sum; // @[MMU.scala 81:29]
  wire  _T_23 = io_smode & _T_22; // @[MMU.scala 81:26]
  wire  uFault = _T_23 & tlb_io_rent_u; // @[MMU.scala 81:37]
  wire  _T_24 = daFault | rFault; // @[MMU.scala 82:25]
  wire  _T_25 = _T_24 | wFault; // @[MMU.scala 82:35]
  wire  vmFault = _T_25 | uFault; // @[MMU.scala 82:55]
  wire  fault = io_en & vmFault; // @[MMU.scala 83:23]
  wire [11:0] voffset = io_vaddr[11:0]; // @[MMU.scala 86:25]
  wire [33:0] _T_27 = {tlb_io_rent_ppn,voffset}; // @[Cat.scala 30:58]
  wire [31:0] tlbAddr = _T_27[31:0]; // @[MMU.scala 87:46]
  wire  _T_28 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_29 = ~tlb_io_valid; // @[MMU.scala 103:28]
  wire  _T_30 = io_lookup & _T_29; // @[MMU.scala 103:25]
  wire [33:0] _T_31 = {io_basePpn, 12'h0}; // @[Paging.scala 41:12]
  wire [11:0] _T_36 = {io_vaddr[31:22], 2'h0}; // @[Paging.scala 41:51]
  wire [33:0] _GEN_82 = {{22'd0}, _T_36}; // @[Paging.scala 41:27]
  wire [33:0] _T_38 = _T_31 + _GEN_82; // @[Paging.scala 41:27]
  wire [33:0] _GEN_1 = _T_30 ? _T_38 : {{2'd0}, addr}; // @[MMU.scala 103:43]
  wire  _GEN_2 = _T_30 | level; // @[MMU.scala 103:43]
  wire [33:0] _GEN_4 = io_en ? _GEN_1 : {{2'd0}, addr}; // @[MMU.scala 101:27]
  wire [33:0] _GEN_7 = io_flush ? {{2'd0}, addr} : _GEN_4; // @[MMU.scala 98:23]
  wire  _T_39 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_40 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_41 = ~pte_v; // @[MMU.scala 118:13]
  wire  _T_42 = ~pte_r; // @[MMU.scala 118:24]
  wire  _T_43 = _T_42 & pte_w; // @[MMU.scala 118:31]
  wire  _T_44 = _T_41 | _T_43; // @[MMU.scala 118:20]
  wire  _T_46 = pte_r | pte_x; // @[MMU.scala 121:26]
  wire  _T_47 = level > 1'h0; // @[MMU.scala 122:21]
  wire  _T_49 = level - 1'h1; // @[MMU.scala 122:58]
  wire [21:0] _T_53 = _T_49 ? pte_ppn : {{12'd0}, pte_ppn[9:0]}; // @[Paging.scala 37:10]
  wire  _T_54 = _T_53 != 22'h0; // @[MMU.scala 122:65]
  wire  _T_55 = _T_47 & _T_54; // @[MMU.scala 122:27]
  wire [21:0] _T_65 = pte_ppn ^ _T_53; // @[Paging.scala 45:12]
  wire [19:0] _T_69 = _T_49 ? io_vaddr[31:12] : {{10'd0}, io_vaddr[21:12]}; // @[Paging.scala 29:10]
  wire [21:0] _GEN_83 = {{2'd0}, _T_69}; // @[Paging.scala 45:40]
  wire [21:0] _T_70 = _T_65 | _GEN_83; // @[Paging.scala 45:40]
  wire  _T_71 = ~level; // @[MMU.scala 134:26]
  wire [33:0] _T_75 = {pte_ppn, 12'h0}; // @[Paging.scala 41:12]
  wire [9:0] _T_79 = _T_49 ? io_vaddr[31:22] : io_vaddr[21:12]; // @[Paging.scala 25:10]
  wire [11:0] _T_80 = {_T_79, 2'h0}; // @[Paging.scala 41:51]
  wire [33:0] _GEN_84 = {{22'd0}, _T_80}; // @[Paging.scala 41:27]
  wire [33:0] _T_82 = _T_75 + _GEN_84; // @[Paging.scala 41:27]
  wire [33:0] _GEN_27 = _T_71 ? {{2'd0}, addr} : _T_82; // @[MMU.scala 134:35]
  wire [33:0] _GEN_37 = _T_46 ? {{2'd0}, addr} : _GEN_27; // @[MMU.scala 121:36]
  wire [33:0] _GEN_47 = _T_44 ? {{2'd0}, addr} : _GEN_37; // @[MMU.scala 118:42]
  wire  _T_85 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_86 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_87 = ~io_flush; // @[MMU.scala 150:13]
  wire [33:0] _GEN_60 = _T_40 ? _GEN_47 : {{2'd0}, addr}; // @[Conditional.scala 39:67]
  wire [33:0] _GEN_70 = _T_39 ? {{2'd0}, addr} : _GEN_60; // @[Conditional.scala 39:67]
  wire [33:0] _GEN_73 = _T_28 ? _GEN_7 : _GEN_70; // @[Conditional.scala 40:58]
  TLB tlb ( // @[MMU.scala 65:19]
    .clock(tlb_clock),
    .reset(tlb_reset),
    .io_flush(tlb_io_flush),
    .io_wen(tlb_io_wen),
    .io_vaddr(tlb_io_vaddr),
    .io_went_ppn(tlb_io_went_ppn),
    .io_went_d(tlb_io_went_d),
    .io_went_a(tlb_io_went_a),
    .io_went_u(tlb_io_went_u),
    .io_went_x(tlb_io_went_x),
    .io_went_w(tlb_io_went_w),
    .io_went_r(tlb_io_went_r),
    .io_valid(tlb_io_valid),
    .io_rent_ppn(tlb_io_rent_ppn),
    .io_rent_d(tlb_io_rent_d),
    .io_rent_a(tlb_io_rent_a),
    .io_rent_u(tlb_io_rent_u),
    .io_rent_x(tlb_io_rent_x),
    .io_rent_w(tlb_io_rent_w),
    .io_rent_r(tlb_io_rent_r)
  );
  assign io_valid = _T_15 | tlbHit; // @[MMU.scala 161:13]
  assign io_fault = valid & fault; // @[MMU.scala 162:13]
  assign io_paddr = io_en ? tlbAddr : io_vaddr; // @[MMU.scala 163:13]
  assign io_data_en = state == 3'h1; // @[MMU.scala 155:17]
  assign io_data_addr = addr; // @[MMU.scala 157:17]
  assign tlb_clock = clock;
  assign tlb_reset = reset;
  assign tlb_io_flush = io_flush; // @[MMU.scala 66:17]
  assign tlb_io_wen = state == 3'h3; // @[MMU.scala 67:17]
  assign tlb_io_vaddr = io_vaddr; // @[MMU.scala 68:17]
  assign tlb_io_went_ppn = entry_ppn; // @[MMU.scala 69:17]
  assign tlb_io_went_d = entry_d; // @[MMU.scala 69:17]
  assign tlb_io_went_a = entry_a; // @[MMU.scala 69:17]
  assign tlb_io_went_u = entry_u; // @[MMU.scala 69:17]
  assign tlb_io_went_x = entry_x; // @[MMU.scala 69:17]
  assign tlb_io_went_w = entry_w; // @[MMU.scala 69:17]
  assign tlb_io_went_r = entry_r; // @[MMU.scala 69:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  entry_ppn = _RAND_1[21:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  entry_d = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  entry_a = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  entry_u = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  entry_x = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  entry_w = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  entry_r = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  addr = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  level = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (_T_28) begin
      if (io_flush) begin
        state <= 3'h4;
      end else if (io_en) begin
        if (_T_30) begin
          state <= 3'h1;
        end
      end
    end else if (_T_39) begin
      if (io_data_valid) begin
        state <= 3'h2;
      end
    end else if (_T_40) begin
      if (_T_44) begin
        state <= 3'h3;
      end else if (_T_46) begin
        state <= 3'h3;
      end else if (_T_71) begin
        state <= 3'h3;
      end else begin
        state <= 3'h1;
      end
    end else if (_T_85) begin
      state <= 3'h0;
    end else if (_T_86) begin
      if (_T_87) begin
        state <= 3'h0;
      end
    end
    if (!(_T_28)) begin
      if (!(_T_39)) begin
        if (_T_40) begin
          if (_T_44) begin
            entry_ppn <= 22'h0;
          end else if (_T_46) begin
            if (_T_55) begin
              entry_ppn <= 22'h0;
            end else if (_T_47) begin
              entry_ppn <= _T_70;
            end else begin
              entry_ppn <= pte_ppn;
            end
          end else if (_T_71) begin
            entry_ppn <= 22'h0;
          end
        end
      end
    end
    if (!(_T_28)) begin
      if (!(_T_39)) begin
        if (_T_40) begin
          if (_T_44) begin
            entry_d <= 1'h0;
          end else if (_T_46) begin
            if (_T_55) begin
              entry_d <= 1'h0;
            end else begin
              entry_d <= pte_d;
            end
          end else if (_T_71) begin
            entry_d <= 1'h0;
          end
        end
      end
    end
    if (!(_T_28)) begin
      if (!(_T_39)) begin
        if (_T_40) begin
          if (_T_44) begin
            entry_a <= 1'h0;
          end else if (_T_46) begin
            if (_T_55) begin
              entry_a <= 1'h0;
            end else begin
              entry_a <= pte_a;
            end
          end else if (_T_71) begin
            entry_a <= 1'h0;
          end
        end
      end
    end
    if (!(_T_28)) begin
      if (!(_T_39)) begin
        if (_T_40) begin
          if (_T_44) begin
            entry_u <= 1'h0;
          end else if (_T_46) begin
            if (_T_55) begin
              entry_u <= 1'h0;
            end else begin
              entry_u <= pte_u;
            end
          end else if (_T_71) begin
            entry_u <= 1'h0;
          end
        end
      end
    end
    if (!(_T_28)) begin
      if (!(_T_39)) begin
        if (_T_40) begin
          if (_T_44) begin
            entry_x <= 1'h0;
          end else if (_T_46) begin
            if (_T_55) begin
              entry_x <= 1'h0;
            end else begin
              entry_x <= pte_x;
            end
          end else if (_T_71) begin
            entry_x <= 1'h0;
          end
        end
      end
    end
    if (!(_T_28)) begin
      if (!(_T_39)) begin
        if (_T_40) begin
          if (_T_44) begin
            entry_w <= 1'h0;
          end else if (_T_46) begin
            if (_T_55) begin
              entry_w <= 1'h0;
            end else begin
              entry_w <= pte_w;
            end
          end else if (_T_71) begin
            entry_w <= 1'h0;
          end
        end
      end
    end
    if (!(_T_28)) begin
      if (!(_T_39)) begin
        if (_T_40) begin
          if (_T_44) begin
            entry_r <= 1'h0;
          end else if (_T_46) begin
            if (_T_55) begin
              entry_r <= 1'h0;
            end else begin
              entry_r <= pte_r;
            end
          end else if (_T_71) begin
            entry_r <= 1'h0;
          end
        end
      end
    end
    addr <= _GEN_73[31:0];
    if (_T_28) begin
      if (!(io_flush)) begin
        if (io_en) begin
          level <= _GEN_2;
        end
      end
    end else if (!(_T_39)) begin
      if (_T_40) begin
        if (!(_T_44)) begin
          if (!(_T_46)) begin
            if (!(_T_71)) begin
              level <= _T_49;
            end
          end
        end
      end
    end
  end
endmodule
module SramMux2(
  input         clock,
  input         io_sel2,
  input         io_in_en,
  output        io_in_valid,
  input  [3:0]  io_in_wen,
  input  [31:0] io_in_addr,
  output [31:0] io_in_rdata,
  input  [31:0] io_in_wdata,
  output        io_out1_en,
  input         io_out1_valid,
  output [3:0]  io_out1_wen,
  output [31:0] io_out1_addr,
  input  [31:0] io_out1_rdata,
  output [31:0] io_out1_wdata,
  output        io_out2_en,
  input         io_out2_valid,
  output [3:0]  io_out2_wen,
  output [31:0] io_out2_addr,
  input  [31:0] io_out2_rdata,
  output [31:0] io_out2_wdata
);
  reg  rdata_sel; // @[SramUtils.scala 16:26]
  reg [31:0] _RAND_0;
  wire  _T_3 = ~io_sel2; // @[SramUtils.scala 22:32]
  assign io_in_valid = io_sel2 ? io_out2_valid : io_out1_valid; // @[SramUtils.scala 18:17]
  assign io_in_rdata = rdata_sel ? io_out2_rdata : io_out1_rdata; // @[SramUtils.scala 20:17]
  assign io_out1_en = io_in_en & _T_3; // @[SramUtils.scala 22:17]
  assign io_out1_wen = io_in_wen; // @[SramUtils.scala 23:17]
  assign io_out1_addr = io_in_addr; // @[SramUtils.scala 24:17]
  assign io_out1_wdata = io_in_wdata; // @[SramUtils.scala 25:17]
  assign io_out2_en = io_in_en & io_sel2; // @[SramUtils.scala 27:17]
  assign io_out2_wen = io_in_wen; // @[SramUtils.scala 28:17]
  assign io_out2_addr = io_in_addr; // @[SramUtils.scala 29:17]
  assign io_out2_wdata = io_in_wdata; // @[SramUtils.scala 30:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rdata_sel = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    rdata_sel <= io_sel2;
  end
endmodule
module BlockMem(
  input         clock,
  input  [3:0]  io_wen,
  input  [10:0] io_addr,
  input  [31:0] io_wdata,
  output [31:0] io_rdata
);
  reg [7:0] mem_0 [0:2047]; // @[BlockMem.scala 20:24]
  reg [31:0] _RAND_0;
  wire [7:0] mem_0__T_11_data; // @[BlockMem.scala 20:24]
  wire [10:0] mem_0__T_11_addr; // @[BlockMem.scala 20:24]
  wire [7:0] mem_0__T_10_data; // @[BlockMem.scala 20:24]
  wire [10:0] mem_0__T_10_addr; // @[BlockMem.scala 20:24]
  wire  mem_0__T_10_mask; // @[BlockMem.scala 20:24]
  wire  mem_0__T_10_en; // @[BlockMem.scala 20:24]
  reg  mem_0__T_11_en_pipe_0;
  reg [31:0] _RAND_1;
  reg [10:0] mem_0__T_11_addr_pipe_0;
  reg [31:0] _RAND_2;
  reg [7:0] mem_1 [0:2047]; // @[BlockMem.scala 20:24]
  reg [31:0] _RAND_3;
  wire [7:0] mem_1__T_11_data; // @[BlockMem.scala 20:24]
  wire [10:0] mem_1__T_11_addr; // @[BlockMem.scala 20:24]
  wire [7:0] mem_1__T_10_data; // @[BlockMem.scala 20:24]
  wire [10:0] mem_1__T_10_addr; // @[BlockMem.scala 20:24]
  wire  mem_1__T_10_mask; // @[BlockMem.scala 20:24]
  wire  mem_1__T_10_en; // @[BlockMem.scala 20:24]
  reg  mem_1__T_11_en_pipe_0;
  reg [31:0] _RAND_4;
  reg [10:0] mem_1__T_11_addr_pipe_0;
  reg [31:0] _RAND_5;
  reg [7:0] mem_2 [0:2047]; // @[BlockMem.scala 20:24]
  reg [31:0] _RAND_6;
  wire [7:0] mem_2__T_11_data; // @[BlockMem.scala 20:24]
  wire [10:0] mem_2__T_11_addr; // @[BlockMem.scala 20:24]
  wire [7:0] mem_2__T_10_data; // @[BlockMem.scala 20:24]
  wire [10:0] mem_2__T_10_addr; // @[BlockMem.scala 20:24]
  wire  mem_2__T_10_mask; // @[BlockMem.scala 20:24]
  wire  mem_2__T_10_en; // @[BlockMem.scala 20:24]
  reg  mem_2__T_11_en_pipe_0;
  reg [31:0] _RAND_7;
  reg [10:0] mem_2__T_11_addr_pipe_0;
  reg [31:0] _RAND_8;
  reg [7:0] mem_3 [0:2047]; // @[BlockMem.scala 20:24]
  reg [31:0] _RAND_9;
  wire [7:0] mem_3__T_11_data; // @[BlockMem.scala 20:24]
  wire [10:0] mem_3__T_11_addr; // @[BlockMem.scala 20:24]
  wire [7:0] mem_3__T_10_data; // @[BlockMem.scala 20:24]
  wire [10:0] mem_3__T_10_addr; // @[BlockMem.scala 20:24]
  wire  mem_3__T_10_mask; // @[BlockMem.scala 20:24]
  wire  mem_3__T_10_en; // @[BlockMem.scala 20:24]
  reg  mem_3__T_11_en_pipe_0;
  reg [31:0] _RAND_10;
  reg [10:0] mem_3__T_11_addr_pipe_0;
  reg [31:0] _RAND_11;
  wire  _T = io_wen != 4'h0; // @[BlockMem.scala 24:18]
  wire [15:0] _T_12 = {mem_1__T_11_data,mem_0__T_11_data}; // @[Cat.scala 30:58]
  wire [15:0] _T_13 = {mem_3__T_11_data,mem_2__T_11_data}; // @[Cat.scala 30:58]
  assign mem_0__T_11_addr = mem_0__T_11_addr_pipe_0;
  assign mem_0__T_11_data = mem_0[mem_0__T_11_addr]; // @[BlockMem.scala 20:24]
  assign mem_0__T_10_data = io_wdata[7:0];
  assign mem_0__T_10_addr = io_addr;
  assign mem_0__T_10_mask = io_wen[0];
  assign mem_0__T_10_en = io_wen != 4'h0;
  assign mem_1__T_11_addr = mem_1__T_11_addr_pipe_0;
  assign mem_1__T_11_data = mem_1[mem_1__T_11_addr]; // @[BlockMem.scala 20:24]
  assign mem_1__T_10_data = io_wdata[15:8];
  assign mem_1__T_10_addr = io_addr;
  assign mem_1__T_10_mask = io_wen[1];
  assign mem_1__T_10_en = io_wen != 4'h0;
  assign mem_2__T_11_addr = mem_2__T_11_addr_pipe_0;
  assign mem_2__T_11_data = mem_2[mem_2__T_11_addr]; // @[BlockMem.scala 20:24]
  assign mem_2__T_10_data = io_wdata[23:16];
  assign mem_2__T_10_addr = io_addr;
  assign mem_2__T_10_mask = io_wen[2];
  assign mem_2__T_10_en = io_wen != 4'h0;
  assign mem_3__T_11_addr = mem_3__T_11_addr_pipe_0;
  assign mem_3__T_11_data = mem_3[mem_3__T_11_addr]; // @[BlockMem.scala 20:24]
  assign mem_3__T_10_data = io_wdata[31:24];
  assign mem_3__T_10_addr = io_addr;
  assign mem_3__T_10_mask = io_wen[3];
  assign mem_3__T_10_en = io_wen != 4'h0;
  assign io_rdata = {_T_13,_T_12}; // @[BlockMem.scala 27:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    mem_0[initvar] = _RAND_0[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem_0__T_11_en_pipe_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  mem_0__T_11_addr_pipe_0 = _RAND_2[10:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    mem_1[initvar] = _RAND_3[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  mem_1__T_11_en_pipe_0 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  mem_1__T_11_addr_pipe_0 = _RAND_5[10:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    mem_2[initvar] = _RAND_6[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  mem_2__T_11_en_pipe_0 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  mem_2__T_11_addr_pipe_0 = _RAND_8[10:0];
  `endif // RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 2048; initvar = initvar+1)
    mem_3[initvar] = _RAND_9[7:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  mem_3__T_11_en_pipe_0 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  mem_3__T_11_addr_pipe_0 = _RAND_11[10:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(mem_0__T_10_en & mem_0__T_10_mask) begin
      mem_0[mem_0__T_10_addr] <= mem_0__T_10_data; // @[BlockMem.scala 20:24]
    end
    if (_T) begin
      mem_0__T_11_en_pipe_0 <= 1'h0;
    end else begin
      mem_0__T_11_en_pipe_0 <= 1'h1;
    end
    if (_T ? 1'h0 : 1'h1) begin
      mem_0__T_11_addr_pipe_0 <= io_addr;
    end
    if(mem_1__T_10_en & mem_1__T_10_mask) begin
      mem_1[mem_1__T_10_addr] <= mem_1__T_10_data; // @[BlockMem.scala 20:24]
    end
    if (_T) begin
      mem_1__T_11_en_pipe_0 <= 1'h0;
    end else begin
      mem_1__T_11_en_pipe_0 <= 1'h1;
    end
    if (_T ? 1'h0 : 1'h1) begin
      mem_1__T_11_addr_pipe_0 <= io_addr;
    end
    if(mem_2__T_10_en & mem_2__T_10_mask) begin
      mem_2[mem_2__T_10_addr] <= mem_2__T_10_data; // @[BlockMem.scala 20:24]
    end
    if (_T) begin
      mem_2__T_11_en_pipe_0 <= 1'h0;
    end else begin
      mem_2__T_11_en_pipe_0 <= 1'h1;
    end
    if (_T ? 1'h0 : 1'h1) begin
      mem_2__T_11_addr_pipe_0 <= io_addr;
    end
    if(mem_3__T_10_en & mem_3__T_10_mask) begin
      mem_3[mem_3__T_10_addr] <= mem_3__T_10_data; // @[BlockMem.scala 20:24]
    end
    if (_T) begin
      mem_3__T_11_en_pipe_0 <= 1'h0;
    end else begin
      mem_3__T_11_en_pipe_0 <= 1'h1;
    end
    if (_T ? 1'h0 : 1'h1) begin
      mem_3__T_11_addr_pipe_0 <= io_addr;
    end
  end
endmodule
module DataCache(
  input         clock,
  input         reset,
  input         io_sram_en,
  output        io_sram_valid,
  input  [3:0]  io_sram_wen,
  input  [31:0] io_sram_addr,
  output [31:0] io_sram_rdata,
  input  [31:0] io_sram_wdata,
  input         io_flush,
  input         io_axi_readAddr_ready,
  output        io_axi_readAddr_valid,
  output [31:0] io_axi_readAddr_bits_addr,
  input         io_axi_readData_valid,
  input  [31:0] io_axi_readData_bits_data,
  input         io_axi_readData_bits_last,
  input         io_axi_writeAddr_ready,
  output        io_axi_writeAddr_valid,
  output [31:0] io_axi_writeAddr_bits_addr,
  input         io_axi_writeData_ready,
  output        io_axi_writeData_valid,
  output [31:0] io_axi_writeData_bits_data,
  output        io_axi_writeData_bits_last
);
  reg [18:0] tag [0:127]; // @[DataCache.scala 39:18]
  reg [31:0] _RAND_0;
  wire [18:0] tag__T_4_data; // @[DataCache.scala 39:18]
  wire [6:0] tag__T_4_addr; // @[DataCache.scala 39:18]
  wire [18:0] tag__T_6_data; // @[DataCache.scala 39:18]
  wire [6:0] tag__T_6_addr; // @[DataCache.scala 39:18]
  wire [18:0] tag__T_261_data; // @[DataCache.scala 39:18]
  wire [6:0] tag__T_261_addr; // @[DataCache.scala 39:18]
  wire [18:0] tag__T_284_data; // @[DataCache.scala 39:18]
  wire [6:0] tag__T_284_addr; // @[DataCache.scala 39:18]
  wire  tag__T_284_mask; // @[DataCache.scala 39:18]
  wire  tag__T_284_en; // @[DataCache.scala 39:18]
  wire  lines_clock; // @[DataCache.scala 40:21]
  wire [3:0] lines_io_wen; // @[DataCache.scala 40:21]
  wire [10:0] lines_io_addr; // @[DataCache.scala 40:21]
  wire [31:0] lines_io_wdata; // @[DataCache.scala 40:21]
  wire [31:0] lines_io_rdata; // @[DataCache.scala 40:21]
  reg [3:0] state; // @[DataCache.scala 34:22]
  reg [31:0] _RAND_1;
  reg  valid_0; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_2;
  reg  valid_1; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_3;
  reg  valid_2; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_4;
  reg  valid_3; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_5;
  reg  valid_4; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_6;
  reg  valid_5; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_7;
  reg  valid_6; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_8;
  reg  valid_7; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_9;
  reg  valid_8; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_10;
  reg  valid_9; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_11;
  reg  valid_10; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_12;
  reg  valid_11; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_13;
  reg  valid_12; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_14;
  reg  valid_13; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_15;
  reg  valid_14; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_16;
  reg  valid_15; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_17;
  reg  valid_16; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_18;
  reg  valid_17; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_19;
  reg  valid_18; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_20;
  reg  valid_19; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_21;
  reg  valid_20; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_22;
  reg  valid_21; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_23;
  reg  valid_22; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_24;
  reg  valid_23; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_25;
  reg  valid_24; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_26;
  reg  valid_25; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_27;
  reg  valid_26; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_28;
  reg  valid_27; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_29;
  reg  valid_28; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_30;
  reg  valid_29; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_31;
  reg  valid_30; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_32;
  reg  valid_31; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_33;
  reg  valid_32; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_34;
  reg  valid_33; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_35;
  reg  valid_34; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_36;
  reg  valid_35; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_37;
  reg  valid_36; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_38;
  reg  valid_37; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_39;
  reg  valid_38; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_40;
  reg  valid_39; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_41;
  reg  valid_40; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_42;
  reg  valid_41; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_43;
  reg  valid_42; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_44;
  reg  valid_43; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_45;
  reg  valid_44; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_46;
  reg  valid_45; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_47;
  reg  valid_46; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_48;
  reg  valid_47; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_49;
  reg  valid_48; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_50;
  reg  valid_49; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_51;
  reg  valid_50; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_52;
  reg  valid_51; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_53;
  reg  valid_52; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_54;
  reg  valid_53; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_55;
  reg  valid_54; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_56;
  reg  valid_55; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_57;
  reg  valid_56; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_58;
  reg  valid_57; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_59;
  reg  valid_58; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_60;
  reg  valid_59; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_61;
  reg  valid_60; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_62;
  reg  valid_61; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_63;
  reg  valid_62; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_64;
  reg  valid_63; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_65;
  reg  valid_64; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_66;
  reg  valid_65; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_67;
  reg  valid_66; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_68;
  reg  valid_67; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_69;
  reg  valid_68; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_70;
  reg  valid_69; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_71;
  reg  valid_70; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_72;
  reg  valid_71; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_73;
  reg  valid_72; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_74;
  reg  valid_73; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_75;
  reg  valid_74; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_76;
  reg  valid_75; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_77;
  reg  valid_76; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_78;
  reg  valid_77; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_79;
  reg  valid_78; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_80;
  reg  valid_79; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_81;
  reg  valid_80; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_82;
  reg  valid_81; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_83;
  reg  valid_82; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_84;
  reg  valid_83; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_85;
  reg  valid_84; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_86;
  reg  valid_85; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_87;
  reg  valid_86; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_88;
  reg  valid_87; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_89;
  reg  valid_88; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_90;
  reg  valid_89; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_91;
  reg  valid_90; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_92;
  reg  valid_91; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_93;
  reg  valid_92; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_94;
  reg  valid_93; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_95;
  reg  valid_94; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_96;
  reg  valid_95; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_97;
  reg  valid_96; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_98;
  reg  valid_97; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_99;
  reg  valid_98; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_100;
  reg  valid_99; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_101;
  reg  valid_100; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_102;
  reg  valid_101; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_103;
  reg  valid_102; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_104;
  reg  valid_103; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_105;
  reg  valid_104; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_106;
  reg  valid_105; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_107;
  reg  valid_106; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_108;
  reg  valid_107; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_109;
  reg  valid_108; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_110;
  reg  valid_109; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_111;
  reg  valid_110; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_112;
  reg  valid_111; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_113;
  reg  valid_112; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_114;
  reg  valid_113; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_115;
  reg  valid_114; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_116;
  reg  valid_115; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_117;
  reg  valid_116; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_118;
  reg  valid_117; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_119;
  reg  valid_118; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_120;
  reg  valid_119; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_121;
  reg  valid_120; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_122;
  reg  valid_121; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_123;
  reg  valid_122; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_124;
  reg  valid_123; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_125;
  reg  valid_124; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_126;
  reg  valid_125; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_127;
  reg  valid_126; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_128;
  reg  valid_127; // @[DataCache.scala 37:22]
  reg [31:0] _RAND_129;
  reg  dirty_0; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_130;
  reg  dirty_1; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_131;
  reg  dirty_2; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_132;
  reg  dirty_3; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_133;
  reg  dirty_4; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_134;
  reg  dirty_5; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_135;
  reg  dirty_6; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_136;
  reg  dirty_7; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_137;
  reg  dirty_8; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_138;
  reg  dirty_9; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_139;
  reg  dirty_10; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_140;
  reg  dirty_11; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_141;
  reg  dirty_12; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_142;
  reg  dirty_13; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_143;
  reg  dirty_14; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_144;
  reg  dirty_15; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_145;
  reg  dirty_16; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_146;
  reg  dirty_17; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_147;
  reg  dirty_18; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_148;
  reg  dirty_19; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_149;
  reg  dirty_20; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_150;
  reg  dirty_21; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_151;
  reg  dirty_22; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_152;
  reg  dirty_23; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_153;
  reg  dirty_24; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_154;
  reg  dirty_25; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_155;
  reg  dirty_26; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_156;
  reg  dirty_27; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_157;
  reg  dirty_28; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_158;
  reg  dirty_29; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_159;
  reg  dirty_30; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_160;
  reg  dirty_31; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_161;
  reg  dirty_32; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_162;
  reg  dirty_33; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_163;
  reg  dirty_34; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_164;
  reg  dirty_35; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_165;
  reg  dirty_36; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_166;
  reg  dirty_37; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_167;
  reg  dirty_38; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_168;
  reg  dirty_39; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_169;
  reg  dirty_40; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_170;
  reg  dirty_41; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_171;
  reg  dirty_42; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_172;
  reg  dirty_43; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_173;
  reg  dirty_44; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_174;
  reg  dirty_45; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_175;
  reg  dirty_46; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_176;
  reg  dirty_47; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_177;
  reg  dirty_48; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_178;
  reg  dirty_49; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_179;
  reg  dirty_50; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_180;
  reg  dirty_51; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_181;
  reg  dirty_52; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_182;
  reg  dirty_53; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_183;
  reg  dirty_54; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_184;
  reg  dirty_55; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_185;
  reg  dirty_56; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_186;
  reg  dirty_57; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_187;
  reg  dirty_58; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_188;
  reg  dirty_59; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_189;
  reg  dirty_60; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_190;
  reg  dirty_61; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_191;
  reg  dirty_62; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_192;
  reg  dirty_63; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_193;
  reg  dirty_64; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_194;
  reg  dirty_65; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_195;
  reg  dirty_66; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_196;
  reg  dirty_67; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_197;
  reg  dirty_68; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_198;
  reg  dirty_69; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_199;
  reg  dirty_70; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_200;
  reg  dirty_71; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_201;
  reg  dirty_72; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_202;
  reg  dirty_73; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_203;
  reg  dirty_74; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_204;
  reg  dirty_75; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_205;
  reg  dirty_76; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_206;
  reg  dirty_77; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_207;
  reg  dirty_78; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_208;
  reg  dirty_79; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_209;
  reg  dirty_80; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_210;
  reg  dirty_81; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_211;
  reg  dirty_82; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_212;
  reg  dirty_83; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_213;
  reg  dirty_84; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_214;
  reg  dirty_85; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_215;
  reg  dirty_86; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_216;
  reg  dirty_87; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_217;
  reg  dirty_88; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_218;
  reg  dirty_89; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_219;
  reg  dirty_90; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_220;
  reg  dirty_91; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_221;
  reg  dirty_92; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_222;
  reg  dirty_93; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_223;
  reg  dirty_94; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_224;
  reg  dirty_95; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_225;
  reg  dirty_96; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_226;
  reg  dirty_97; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_227;
  reg  dirty_98; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_228;
  reg  dirty_99; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_229;
  reg  dirty_100; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_230;
  reg  dirty_101; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_231;
  reg  dirty_102; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_232;
  reg  dirty_103; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_233;
  reg  dirty_104; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_234;
  reg  dirty_105; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_235;
  reg  dirty_106; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_236;
  reg  dirty_107; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_237;
  reg  dirty_108; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_238;
  reg  dirty_109; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_239;
  reg  dirty_110; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_240;
  reg  dirty_111; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_241;
  reg  dirty_112; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_242;
  reg  dirty_113; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_243;
  reg  dirty_114; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_244;
  reg  dirty_115; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_245;
  reg  dirty_116; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_246;
  reg  dirty_117; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_247;
  reg  dirty_118; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_248;
  reg  dirty_119; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_249;
  reg  dirty_120; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_250;
  reg  dirty_121; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_251;
  reg  dirty_122; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_252;
  reg  dirty_123; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_253;
  reg  dirty_124; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_254;
  reg  dirty_125; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_255;
  reg  dirty_126; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_256;
  reg  dirty_127; // @[DataCache.scala 38:18]
  reg [31:0] _RAND_257;
  reg [4:0] dataOffset; // @[DataCache.scala 43:24]
  reg [31:0] _RAND_258;
  reg [4:0] lastOffset; // @[DataCache.scala 44:24]
  reg [31:0] _RAND_259;
  wire [3:0] dataOfsRef = dataOffset[3:0]; // @[DataCache.scala 45:31]
  reg  aren; // @[DataCache.scala 46:28]
  reg [31:0] _RAND_260;
  reg [31:0] raddr; // @[DataCache.scala 47:24]
  reg [31:0] _RAND_261;
  reg  awen; // @[DataCache.scala 48:28]
  reg [31:0] _RAND_262;
  reg [31:0] waddr; // @[DataCache.scala 49:24]
  reg [31:0] _RAND_263;
  reg  wen; // @[DataCache.scala 50:28]
  reg [31:0] _RAND_264;
  wire  _T_1 = dataOffset == 5'h10; // @[DataCache.scala 51:39]
  wire  wlast = wen & _T_1; // @[DataCache.scala 51:25]
  reg [31:0] sramAddr; // @[DataCache.scala 54:24]
  reg [31:0] _RAND_265;
  wire  _T_2 = state == 4'h0; // @[DataCache.scala 55:31]
  wire [31:0] selAddr = _T_2 ? io_sram_addr : sramAddr; // @[DataCache.scala 55:24]
  wire [18:0] tagSel = selAddr[31:13]; // @[DataCache.scala 56:28]
  wire [6:0] lineSel = selAddr[12:6]; // @[DataCache.scala 58:28]
  wire [10:0] lineDataSel = selAddr[12:2]; // @[DataCache.scala 60:28]
  wire [10:0] dataSel = {lineSel,dataOfsRef}; // @[Cat.scala 30:58]
  wire [31:0] startRaddr = {tagSel,lineSel,6'h0}; // @[Cat.scala 30:58]
  wire [31:0] startWaddr = {tag__T_4_data,lineSel,6'h0}; // @[Cat.scala 30:58]
  wire  _T_7 = tag__T_6_data == tagSel; // @[DataCache.scala 67:50]
  wire  _GEN_1 = 7'h1 == lineSel ? valid_1 : valid_0; // @[DataCache.scala 67:34]
  wire  _GEN_2 = 7'h2 == lineSel ? valid_2 : _GEN_1; // @[DataCache.scala 67:34]
  wire  _GEN_3 = 7'h3 == lineSel ? valid_3 : _GEN_2; // @[DataCache.scala 67:34]
  wire  _GEN_4 = 7'h4 == lineSel ? valid_4 : _GEN_3; // @[DataCache.scala 67:34]
  wire  _GEN_5 = 7'h5 == lineSel ? valid_5 : _GEN_4; // @[DataCache.scala 67:34]
  wire  _GEN_6 = 7'h6 == lineSel ? valid_6 : _GEN_5; // @[DataCache.scala 67:34]
  wire  _GEN_7 = 7'h7 == lineSel ? valid_7 : _GEN_6; // @[DataCache.scala 67:34]
  wire  _GEN_8 = 7'h8 == lineSel ? valid_8 : _GEN_7; // @[DataCache.scala 67:34]
  wire  _GEN_9 = 7'h9 == lineSel ? valid_9 : _GEN_8; // @[DataCache.scala 67:34]
  wire  _GEN_10 = 7'ha == lineSel ? valid_10 : _GEN_9; // @[DataCache.scala 67:34]
  wire  _GEN_11 = 7'hb == lineSel ? valid_11 : _GEN_10; // @[DataCache.scala 67:34]
  wire  _GEN_12 = 7'hc == lineSel ? valid_12 : _GEN_11; // @[DataCache.scala 67:34]
  wire  _GEN_13 = 7'hd == lineSel ? valid_13 : _GEN_12; // @[DataCache.scala 67:34]
  wire  _GEN_14 = 7'he == lineSel ? valid_14 : _GEN_13; // @[DataCache.scala 67:34]
  wire  _GEN_15 = 7'hf == lineSel ? valid_15 : _GEN_14; // @[DataCache.scala 67:34]
  wire  _GEN_16 = 7'h10 == lineSel ? valid_16 : _GEN_15; // @[DataCache.scala 67:34]
  wire  _GEN_17 = 7'h11 == lineSel ? valid_17 : _GEN_16; // @[DataCache.scala 67:34]
  wire  _GEN_18 = 7'h12 == lineSel ? valid_18 : _GEN_17; // @[DataCache.scala 67:34]
  wire  _GEN_19 = 7'h13 == lineSel ? valid_19 : _GEN_18; // @[DataCache.scala 67:34]
  wire  _GEN_20 = 7'h14 == lineSel ? valid_20 : _GEN_19; // @[DataCache.scala 67:34]
  wire  _GEN_21 = 7'h15 == lineSel ? valid_21 : _GEN_20; // @[DataCache.scala 67:34]
  wire  _GEN_22 = 7'h16 == lineSel ? valid_22 : _GEN_21; // @[DataCache.scala 67:34]
  wire  _GEN_23 = 7'h17 == lineSel ? valid_23 : _GEN_22; // @[DataCache.scala 67:34]
  wire  _GEN_24 = 7'h18 == lineSel ? valid_24 : _GEN_23; // @[DataCache.scala 67:34]
  wire  _GEN_25 = 7'h19 == lineSel ? valid_25 : _GEN_24; // @[DataCache.scala 67:34]
  wire  _GEN_26 = 7'h1a == lineSel ? valid_26 : _GEN_25; // @[DataCache.scala 67:34]
  wire  _GEN_27 = 7'h1b == lineSel ? valid_27 : _GEN_26; // @[DataCache.scala 67:34]
  wire  _GEN_28 = 7'h1c == lineSel ? valid_28 : _GEN_27; // @[DataCache.scala 67:34]
  wire  _GEN_29 = 7'h1d == lineSel ? valid_29 : _GEN_28; // @[DataCache.scala 67:34]
  wire  _GEN_30 = 7'h1e == lineSel ? valid_30 : _GEN_29; // @[DataCache.scala 67:34]
  wire  _GEN_31 = 7'h1f == lineSel ? valid_31 : _GEN_30; // @[DataCache.scala 67:34]
  wire  _GEN_32 = 7'h20 == lineSel ? valid_32 : _GEN_31; // @[DataCache.scala 67:34]
  wire  _GEN_33 = 7'h21 == lineSel ? valid_33 : _GEN_32; // @[DataCache.scala 67:34]
  wire  _GEN_34 = 7'h22 == lineSel ? valid_34 : _GEN_33; // @[DataCache.scala 67:34]
  wire  _GEN_35 = 7'h23 == lineSel ? valid_35 : _GEN_34; // @[DataCache.scala 67:34]
  wire  _GEN_36 = 7'h24 == lineSel ? valid_36 : _GEN_35; // @[DataCache.scala 67:34]
  wire  _GEN_37 = 7'h25 == lineSel ? valid_37 : _GEN_36; // @[DataCache.scala 67:34]
  wire  _GEN_38 = 7'h26 == lineSel ? valid_38 : _GEN_37; // @[DataCache.scala 67:34]
  wire  _GEN_39 = 7'h27 == lineSel ? valid_39 : _GEN_38; // @[DataCache.scala 67:34]
  wire  _GEN_40 = 7'h28 == lineSel ? valid_40 : _GEN_39; // @[DataCache.scala 67:34]
  wire  _GEN_41 = 7'h29 == lineSel ? valid_41 : _GEN_40; // @[DataCache.scala 67:34]
  wire  _GEN_42 = 7'h2a == lineSel ? valid_42 : _GEN_41; // @[DataCache.scala 67:34]
  wire  _GEN_43 = 7'h2b == lineSel ? valid_43 : _GEN_42; // @[DataCache.scala 67:34]
  wire  _GEN_44 = 7'h2c == lineSel ? valid_44 : _GEN_43; // @[DataCache.scala 67:34]
  wire  _GEN_45 = 7'h2d == lineSel ? valid_45 : _GEN_44; // @[DataCache.scala 67:34]
  wire  _GEN_46 = 7'h2e == lineSel ? valid_46 : _GEN_45; // @[DataCache.scala 67:34]
  wire  _GEN_47 = 7'h2f == lineSel ? valid_47 : _GEN_46; // @[DataCache.scala 67:34]
  wire  _GEN_48 = 7'h30 == lineSel ? valid_48 : _GEN_47; // @[DataCache.scala 67:34]
  wire  _GEN_49 = 7'h31 == lineSel ? valid_49 : _GEN_48; // @[DataCache.scala 67:34]
  wire  _GEN_50 = 7'h32 == lineSel ? valid_50 : _GEN_49; // @[DataCache.scala 67:34]
  wire  _GEN_51 = 7'h33 == lineSel ? valid_51 : _GEN_50; // @[DataCache.scala 67:34]
  wire  _GEN_52 = 7'h34 == lineSel ? valid_52 : _GEN_51; // @[DataCache.scala 67:34]
  wire  _GEN_53 = 7'h35 == lineSel ? valid_53 : _GEN_52; // @[DataCache.scala 67:34]
  wire  _GEN_54 = 7'h36 == lineSel ? valid_54 : _GEN_53; // @[DataCache.scala 67:34]
  wire  _GEN_55 = 7'h37 == lineSel ? valid_55 : _GEN_54; // @[DataCache.scala 67:34]
  wire  _GEN_56 = 7'h38 == lineSel ? valid_56 : _GEN_55; // @[DataCache.scala 67:34]
  wire  _GEN_57 = 7'h39 == lineSel ? valid_57 : _GEN_56; // @[DataCache.scala 67:34]
  wire  _GEN_58 = 7'h3a == lineSel ? valid_58 : _GEN_57; // @[DataCache.scala 67:34]
  wire  _GEN_59 = 7'h3b == lineSel ? valid_59 : _GEN_58; // @[DataCache.scala 67:34]
  wire  _GEN_60 = 7'h3c == lineSel ? valid_60 : _GEN_59; // @[DataCache.scala 67:34]
  wire  _GEN_61 = 7'h3d == lineSel ? valid_61 : _GEN_60; // @[DataCache.scala 67:34]
  wire  _GEN_62 = 7'h3e == lineSel ? valid_62 : _GEN_61; // @[DataCache.scala 67:34]
  wire  _GEN_63 = 7'h3f == lineSel ? valid_63 : _GEN_62; // @[DataCache.scala 67:34]
  wire  _GEN_64 = 7'h40 == lineSel ? valid_64 : _GEN_63; // @[DataCache.scala 67:34]
  wire  _GEN_65 = 7'h41 == lineSel ? valid_65 : _GEN_64; // @[DataCache.scala 67:34]
  wire  _GEN_66 = 7'h42 == lineSel ? valid_66 : _GEN_65; // @[DataCache.scala 67:34]
  wire  _GEN_67 = 7'h43 == lineSel ? valid_67 : _GEN_66; // @[DataCache.scala 67:34]
  wire  _GEN_68 = 7'h44 == lineSel ? valid_68 : _GEN_67; // @[DataCache.scala 67:34]
  wire  _GEN_69 = 7'h45 == lineSel ? valid_69 : _GEN_68; // @[DataCache.scala 67:34]
  wire  _GEN_70 = 7'h46 == lineSel ? valid_70 : _GEN_69; // @[DataCache.scala 67:34]
  wire  _GEN_71 = 7'h47 == lineSel ? valid_71 : _GEN_70; // @[DataCache.scala 67:34]
  wire  _GEN_72 = 7'h48 == lineSel ? valid_72 : _GEN_71; // @[DataCache.scala 67:34]
  wire  _GEN_73 = 7'h49 == lineSel ? valid_73 : _GEN_72; // @[DataCache.scala 67:34]
  wire  _GEN_74 = 7'h4a == lineSel ? valid_74 : _GEN_73; // @[DataCache.scala 67:34]
  wire  _GEN_75 = 7'h4b == lineSel ? valid_75 : _GEN_74; // @[DataCache.scala 67:34]
  wire  _GEN_76 = 7'h4c == lineSel ? valid_76 : _GEN_75; // @[DataCache.scala 67:34]
  wire  _GEN_77 = 7'h4d == lineSel ? valid_77 : _GEN_76; // @[DataCache.scala 67:34]
  wire  _GEN_78 = 7'h4e == lineSel ? valid_78 : _GEN_77; // @[DataCache.scala 67:34]
  wire  _GEN_79 = 7'h4f == lineSel ? valid_79 : _GEN_78; // @[DataCache.scala 67:34]
  wire  _GEN_80 = 7'h50 == lineSel ? valid_80 : _GEN_79; // @[DataCache.scala 67:34]
  wire  _GEN_81 = 7'h51 == lineSel ? valid_81 : _GEN_80; // @[DataCache.scala 67:34]
  wire  _GEN_82 = 7'h52 == lineSel ? valid_82 : _GEN_81; // @[DataCache.scala 67:34]
  wire  _GEN_83 = 7'h53 == lineSel ? valid_83 : _GEN_82; // @[DataCache.scala 67:34]
  wire  _GEN_84 = 7'h54 == lineSel ? valid_84 : _GEN_83; // @[DataCache.scala 67:34]
  wire  _GEN_85 = 7'h55 == lineSel ? valid_85 : _GEN_84; // @[DataCache.scala 67:34]
  wire  _GEN_86 = 7'h56 == lineSel ? valid_86 : _GEN_85; // @[DataCache.scala 67:34]
  wire  _GEN_87 = 7'h57 == lineSel ? valid_87 : _GEN_86; // @[DataCache.scala 67:34]
  wire  _GEN_88 = 7'h58 == lineSel ? valid_88 : _GEN_87; // @[DataCache.scala 67:34]
  wire  _GEN_89 = 7'h59 == lineSel ? valid_89 : _GEN_88; // @[DataCache.scala 67:34]
  wire  _GEN_90 = 7'h5a == lineSel ? valid_90 : _GEN_89; // @[DataCache.scala 67:34]
  wire  _GEN_91 = 7'h5b == lineSel ? valid_91 : _GEN_90; // @[DataCache.scala 67:34]
  wire  _GEN_92 = 7'h5c == lineSel ? valid_92 : _GEN_91; // @[DataCache.scala 67:34]
  wire  _GEN_93 = 7'h5d == lineSel ? valid_93 : _GEN_92; // @[DataCache.scala 67:34]
  wire  _GEN_94 = 7'h5e == lineSel ? valid_94 : _GEN_93; // @[DataCache.scala 67:34]
  wire  _GEN_95 = 7'h5f == lineSel ? valid_95 : _GEN_94; // @[DataCache.scala 67:34]
  wire  _GEN_96 = 7'h60 == lineSel ? valid_96 : _GEN_95; // @[DataCache.scala 67:34]
  wire  _GEN_97 = 7'h61 == lineSel ? valid_97 : _GEN_96; // @[DataCache.scala 67:34]
  wire  _GEN_98 = 7'h62 == lineSel ? valid_98 : _GEN_97; // @[DataCache.scala 67:34]
  wire  _GEN_99 = 7'h63 == lineSel ? valid_99 : _GEN_98; // @[DataCache.scala 67:34]
  wire  _GEN_100 = 7'h64 == lineSel ? valid_100 : _GEN_99; // @[DataCache.scala 67:34]
  wire  _GEN_101 = 7'h65 == lineSel ? valid_101 : _GEN_100; // @[DataCache.scala 67:34]
  wire  _GEN_102 = 7'h66 == lineSel ? valid_102 : _GEN_101; // @[DataCache.scala 67:34]
  wire  _GEN_103 = 7'h67 == lineSel ? valid_103 : _GEN_102; // @[DataCache.scala 67:34]
  wire  _GEN_104 = 7'h68 == lineSel ? valid_104 : _GEN_103; // @[DataCache.scala 67:34]
  wire  _GEN_105 = 7'h69 == lineSel ? valid_105 : _GEN_104; // @[DataCache.scala 67:34]
  wire  _GEN_106 = 7'h6a == lineSel ? valid_106 : _GEN_105; // @[DataCache.scala 67:34]
  wire  _GEN_107 = 7'h6b == lineSel ? valid_107 : _GEN_106; // @[DataCache.scala 67:34]
  wire  _GEN_108 = 7'h6c == lineSel ? valid_108 : _GEN_107; // @[DataCache.scala 67:34]
  wire  _GEN_109 = 7'h6d == lineSel ? valid_109 : _GEN_108; // @[DataCache.scala 67:34]
  wire  _GEN_110 = 7'h6e == lineSel ? valid_110 : _GEN_109; // @[DataCache.scala 67:34]
  wire  _GEN_111 = 7'h6f == lineSel ? valid_111 : _GEN_110; // @[DataCache.scala 67:34]
  wire  _GEN_112 = 7'h70 == lineSel ? valid_112 : _GEN_111; // @[DataCache.scala 67:34]
  wire  _GEN_113 = 7'h71 == lineSel ? valid_113 : _GEN_112; // @[DataCache.scala 67:34]
  wire  _GEN_114 = 7'h72 == lineSel ? valid_114 : _GEN_113; // @[DataCache.scala 67:34]
  wire  _GEN_115 = 7'h73 == lineSel ? valid_115 : _GEN_114; // @[DataCache.scala 67:34]
  wire  _GEN_116 = 7'h74 == lineSel ? valid_116 : _GEN_115; // @[DataCache.scala 67:34]
  wire  _GEN_117 = 7'h75 == lineSel ? valid_117 : _GEN_116; // @[DataCache.scala 67:34]
  wire  _GEN_118 = 7'h76 == lineSel ? valid_118 : _GEN_117; // @[DataCache.scala 67:34]
  wire  _GEN_119 = 7'h77 == lineSel ? valid_119 : _GEN_118; // @[DataCache.scala 67:34]
  wire  _GEN_120 = 7'h78 == lineSel ? valid_120 : _GEN_119; // @[DataCache.scala 67:34]
  wire  _GEN_121 = 7'h79 == lineSel ? valid_121 : _GEN_120; // @[DataCache.scala 67:34]
  wire  _GEN_122 = 7'h7a == lineSel ? valid_122 : _GEN_121; // @[DataCache.scala 67:34]
  wire  _GEN_123 = 7'h7b == lineSel ? valid_123 : _GEN_122; // @[DataCache.scala 67:34]
  wire  _GEN_124 = 7'h7c == lineSel ? valid_124 : _GEN_123; // @[DataCache.scala 67:34]
  wire  _GEN_125 = 7'h7d == lineSel ? valid_125 : _GEN_124; // @[DataCache.scala 67:34]
  wire  _GEN_126 = 7'h7e == lineSel ? valid_126 : _GEN_125; // @[DataCache.scala 67:34]
  wire  _GEN_127 = 7'h7f == lineSel ? valid_127 : _GEN_126; // @[DataCache.scala 67:34]
  wire  cacheHit = _GEN_127 & _T_7; // @[DataCache.scala 67:34]
  wire  realDirty_0 = valid_0 & dirty_0; // @[DataCache.scala 68:59]
  wire  realDirty_1 = valid_1 & dirty_1; // @[DataCache.scala 68:59]
  wire  realDirty_2 = valid_2 & dirty_2; // @[DataCache.scala 68:59]
  wire  realDirty_3 = valid_3 & dirty_3; // @[DataCache.scala 68:59]
  wire  realDirty_4 = valid_4 & dirty_4; // @[DataCache.scala 68:59]
  wire  realDirty_5 = valid_5 & dirty_5; // @[DataCache.scala 68:59]
  wire  realDirty_6 = valid_6 & dirty_6; // @[DataCache.scala 68:59]
  wire  realDirty_7 = valid_7 & dirty_7; // @[DataCache.scala 68:59]
  wire  realDirty_8 = valid_8 & dirty_8; // @[DataCache.scala 68:59]
  wire  realDirty_9 = valid_9 & dirty_9; // @[DataCache.scala 68:59]
  wire  realDirty_10 = valid_10 & dirty_10; // @[DataCache.scala 68:59]
  wire  realDirty_11 = valid_11 & dirty_11; // @[DataCache.scala 68:59]
  wire  realDirty_12 = valid_12 & dirty_12; // @[DataCache.scala 68:59]
  wire  realDirty_13 = valid_13 & dirty_13; // @[DataCache.scala 68:59]
  wire  realDirty_14 = valid_14 & dirty_14; // @[DataCache.scala 68:59]
  wire  realDirty_15 = valid_15 & dirty_15; // @[DataCache.scala 68:59]
  wire  realDirty_16 = valid_16 & dirty_16; // @[DataCache.scala 68:59]
  wire  realDirty_17 = valid_17 & dirty_17; // @[DataCache.scala 68:59]
  wire  realDirty_18 = valid_18 & dirty_18; // @[DataCache.scala 68:59]
  wire  realDirty_19 = valid_19 & dirty_19; // @[DataCache.scala 68:59]
  wire  realDirty_20 = valid_20 & dirty_20; // @[DataCache.scala 68:59]
  wire  realDirty_21 = valid_21 & dirty_21; // @[DataCache.scala 68:59]
  wire  realDirty_22 = valid_22 & dirty_22; // @[DataCache.scala 68:59]
  wire  realDirty_23 = valid_23 & dirty_23; // @[DataCache.scala 68:59]
  wire  realDirty_24 = valid_24 & dirty_24; // @[DataCache.scala 68:59]
  wire  realDirty_25 = valid_25 & dirty_25; // @[DataCache.scala 68:59]
  wire  realDirty_26 = valid_26 & dirty_26; // @[DataCache.scala 68:59]
  wire  realDirty_27 = valid_27 & dirty_27; // @[DataCache.scala 68:59]
  wire  realDirty_28 = valid_28 & dirty_28; // @[DataCache.scala 68:59]
  wire  realDirty_29 = valid_29 & dirty_29; // @[DataCache.scala 68:59]
  wire  realDirty_30 = valid_30 & dirty_30; // @[DataCache.scala 68:59]
  wire  realDirty_31 = valid_31 & dirty_31; // @[DataCache.scala 68:59]
  wire  realDirty_32 = valid_32 & dirty_32; // @[DataCache.scala 68:59]
  wire  realDirty_33 = valid_33 & dirty_33; // @[DataCache.scala 68:59]
  wire  realDirty_34 = valid_34 & dirty_34; // @[DataCache.scala 68:59]
  wire  realDirty_35 = valid_35 & dirty_35; // @[DataCache.scala 68:59]
  wire  realDirty_36 = valid_36 & dirty_36; // @[DataCache.scala 68:59]
  wire  realDirty_37 = valid_37 & dirty_37; // @[DataCache.scala 68:59]
  wire  realDirty_38 = valid_38 & dirty_38; // @[DataCache.scala 68:59]
  wire  realDirty_39 = valid_39 & dirty_39; // @[DataCache.scala 68:59]
  wire  realDirty_40 = valid_40 & dirty_40; // @[DataCache.scala 68:59]
  wire  realDirty_41 = valid_41 & dirty_41; // @[DataCache.scala 68:59]
  wire  realDirty_42 = valid_42 & dirty_42; // @[DataCache.scala 68:59]
  wire  realDirty_43 = valid_43 & dirty_43; // @[DataCache.scala 68:59]
  wire  realDirty_44 = valid_44 & dirty_44; // @[DataCache.scala 68:59]
  wire  realDirty_45 = valid_45 & dirty_45; // @[DataCache.scala 68:59]
  wire  realDirty_46 = valid_46 & dirty_46; // @[DataCache.scala 68:59]
  wire  realDirty_47 = valid_47 & dirty_47; // @[DataCache.scala 68:59]
  wire  realDirty_48 = valid_48 & dirty_48; // @[DataCache.scala 68:59]
  wire  realDirty_49 = valid_49 & dirty_49; // @[DataCache.scala 68:59]
  wire  realDirty_50 = valid_50 & dirty_50; // @[DataCache.scala 68:59]
  wire  realDirty_51 = valid_51 & dirty_51; // @[DataCache.scala 68:59]
  wire  realDirty_52 = valid_52 & dirty_52; // @[DataCache.scala 68:59]
  wire  realDirty_53 = valid_53 & dirty_53; // @[DataCache.scala 68:59]
  wire  realDirty_54 = valid_54 & dirty_54; // @[DataCache.scala 68:59]
  wire  realDirty_55 = valid_55 & dirty_55; // @[DataCache.scala 68:59]
  wire  realDirty_56 = valid_56 & dirty_56; // @[DataCache.scala 68:59]
  wire  realDirty_57 = valid_57 & dirty_57; // @[DataCache.scala 68:59]
  wire  realDirty_58 = valid_58 & dirty_58; // @[DataCache.scala 68:59]
  wire  realDirty_59 = valid_59 & dirty_59; // @[DataCache.scala 68:59]
  wire  realDirty_60 = valid_60 & dirty_60; // @[DataCache.scala 68:59]
  wire  realDirty_61 = valid_61 & dirty_61; // @[DataCache.scala 68:59]
  wire  realDirty_62 = valid_62 & dirty_62; // @[DataCache.scala 68:59]
  wire  realDirty_63 = valid_63 & dirty_63; // @[DataCache.scala 68:59]
  wire  realDirty_64 = valid_64 & dirty_64; // @[DataCache.scala 68:59]
  wire  realDirty_65 = valid_65 & dirty_65; // @[DataCache.scala 68:59]
  wire  realDirty_66 = valid_66 & dirty_66; // @[DataCache.scala 68:59]
  wire  realDirty_67 = valid_67 & dirty_67; // @[DataCache.scala 68:59]
  wire  realDirty_68 = valid_68 & dirty_68; // @[DataCache.scala 68:59]
  wire  realDirty_69 = valid_69 & dirty_69; // @[DataCache.scala 68:59]
  wire  realDirty_70 = valid_70 & dirty_70; // @[DataCache.scala 68:59]
  wire  realDirty_71 = valid_71 & dirty_71; // @[DataCache.scala 68:59]
  wire  realDirty_72 = valid_72 & dirty_72; // @[DataCache.scala 68:59]
  wire  realDirty_73 = valid_73 & dirty_73; // @[DataCache.scala 68:59]
  wire  realDirty_74 = valid_74 & dirty_74; // @[DataCache.scala 68:59]
  wire  realDirty_75 = valid_75 & dirty_75; // @[DataCache.scala 68:59]
  wire  realDirty_76 = valid_76 & dirty_76; // @[DataCache.scala 68:59]
  wire  realDirty_77 = valid_77 & dirty_77; // @[DataCache.scala 68:59]
  wire  realDirty_78 = valid_78 & dirty_78; // @[DataCache.scala 68:59]
  wire  realDirty_79 = valid_79 & dirty_79; // @[DataCache.scala 68:59]
  wire  realDirty_80 = valid_80 & dirty_80; // @[DataCache.scala 68:59]
  wire  realDirty_81 = valid_81 & dirty_81; // @[DataCache.scala 68:59]
  wire  realDirty_82 = valid_82 & dirty_82; // @[DataCache.scala 68:59]
  wire  realDirty_83 = valid_83 & dirty_83; // @[DataCache.scala 68:59]
  wire  realDirty_84 = valid_84 & dirty_84; // @[DataCache.scala 68:59]
  wire  realDirty_85 = valid_85 & dirty_85; // @[DataCache.scala 68:59]
  wire  realDirty_86 = valid_86 & dirty_86; // @[DataCache.scala 68:59]
  wire  realDirty_87 = valid_87 & dirty_87; // @[DataCache.scala 68:59]
  wire  realDirty_88 = valid_88 & dirty_88; // @[DataCache.scala 68:59]
  wire  realDirty_89 = valid_89 & dirty_89; // @[DataCache.scala 68:59]
  wire  realDirty_90 = valid_90 & dirty_90; // @[DataCache.scala 68:59]
  wire  realDirty_91 = valid_91 & dirty_91; // @[DataCache.scala 68:59]
  wire  realDirty_92 = valid_92 & dirty_92; // @[DataCache.scala 68:59]
  wire  realDirty_93 = valid_93 & dirty_93; // @[DataCache.scala 68:59]
  wire  realDirty_94 = valid_94 & dirty_94; // @[DataCache.scala 68:59]
  wire  realDirty_95 = valid_95 & dirty_95; // @[DataCache.scala 68:59]
  wire  realDirty_96 = valid_96 & dirty_96; // @[DataCache.scala 68:59]
  wire  realDirty_97 = valid_97 & dirty_97; // @[DataCache.scala 68:59]
  wire  realDirty_98 = valid_98 & dirty_98; // @[DataCache.scala 68:59]
  wire  realDirty_99 = valid_99 & dirty_99; // @[DataCache.scala 68:59]
  wire  realDirty_100 = valid_100 & dirty_100; // @[DataCache.scala 68:59]
  wire  realDirty_101 = valid_101 & dirty_101; // @[DataCache.scala 68:59]
  wire  realDirty_102 = valid_102 & dirty_102; // @[DataCache.scala 68:59]
  wire  realDirty_103 = valid_103 & dirty_103; // @[DataCache.scala 68:59]
  wire  realDirty_104 = valid_104 & dirty_104; // @[DataCache.scala 68:59]
  wire  realDirty_105 = valid_105 & dirty_105; // @[DataCache.scala 68:59]
  wire  realDirty_106 = valid_106 & dirty_106; // @[DataCache.scala 68:59]
  wire  realDirty_107 = valid_107 & dirty_107; // @[DataCache.scala 68:59]
  wire  realDirty_108 = valid_108 & dirty_108; // @[DataCache.scala 68:59]
  wire  realDirty_109 = valid_109 & dirty_109; // @[DataCache.scala 68:59]
  wire  realDirty_110 = valid_110 & dirty_110; // @[DataCache.scala 68:59]
  wire  realDirty_111 = valid_111 & dirty_111; // @[DataCache.scala 68:59]
  wire  realDirty_112 = valid_112 & dirty_112; // @[DataCache.scala 68:59]
  wire  realDirty_113 = valid_113 & dirty_113; // @[DataCache.scala 68:59]
  wire  realDirty_114 = valid_114 & dirty_114; // @[DataCache.scala 68:59]
  wire  realDirty_115 = valid_115 & dirty_115; // @[DataCache.scala 68:59]
  wire  realDirty_116 = valid_116 & dirty_116; // @[DataCache.scala 68:59]
  wire  realDirty_117 = valid_117 & dirty_117; // @[DataCache.scala 68:59]
  wire  realDirty_118 = valid_118 & dirty_118; // @[DataCache.scala 68:59]
  wire  realDirty_119 = valid_119 & dirty_119; // @[DataCache.scala 68:59]
  wire  realDirty_120 = valid_120 & dirty_120; // @[DataCache.scala 68:59]
  wire  realDirty_121 = valid_121 & dirty_121; // @[DataCache.scala 68:59]
  wire  realDirty_122 = valid_122 & dirty_122; // @[DataCache.scala 68:59]
  wire  realDirty_123 = valid_123 & dirty_123; // @[DataCache.scala 68:59]
  wire  realDirty_124 = valid_124 & dirty_124; // @[DataCache.scala 68:59]
  wire  realDirty_125 = valid_125 & dirty_125; // @[DataCache.scala 68:59]
  wire  realDirty_126 = valid_126 & dirty_126; // @[DataCache.scala 68:59]
  wire  realDirty_127 = valid_127 & dirty_127; // @[DataCache.scala 68:59]
  wire  _T_8 = realDirty_0 | realDirty_1; // @[DataCache.scala 69:37]
  wire  _T_9 = _T_8 | realDirty_2; // @[DataCache.scala 69:37]
  wire  _T_10 = _T_9 | realDirty_3; // @[DataCache.scala 69:37]
  wire  _T_11 = _T_10 | realDirty_4; // @[DataCache.scala 69:37]
  wire  _T_12 = _T_11 | realDirty_5; // @[DataCache.scala 69:37]
  wire  _T_13 = _T_12 | realDirty_6; // @[DataCache.scala 69:37]
  wire  _T_14 = _T_13 | realDirty_7; // @[DataCache.scala 69:37]
  wire  _T_15 = _T_14 | realDirty_8; // @[DataCache.scala 69:37]
  wire  _T_16 = _T_15 | realDirty_9; // @[DataCache.scala 69:37]
  wire  _T_17 = _T_16 | realDirty_10; // @[DataCache.scala 69:37]
  wire  _T_18 = _T_17 | realDirty_11; // @[DataCache.scala 69:37]
  wire  _T_19 = _T_18 | realDirty_12; // @[DataCache.scala 69:37]
  wire  _T_20 = _T_19 | realDirty_13; // @[DataCache.scala 69:37]
  wire  _T_21 = _T_20 | realDirty_14; // @[DataCache.scala 69:37]
  wire  _T_22 = _T_21 | realDirty_15; // @[DataCache.scala 69:37]
  wire  _T_23 = _T_22 | realDirty_16; // @[DataCache.scala 69:37]
  wire  _T_24 = _T_23 | realDirty_17; // @[DataCache.scala 69:37]
  wire  _T_25 = _T_24 | realDirty_18; // @[DataCache.scala 69:37]
  wire  _T_26 = _T_25 | realDirty_19; // @[DataCache.scala 69:37]
  wire  _T_27 = _T_26 | realDirty_20; // @[DataCache.scala 69:37]
  wire  _T_28 = _T_27 | realDirty_21; // @[DataCache.scala 69:37]
  wire  _T_29 = _T_28 | realDirty_22; // @[DataCache.scala 69:37]
  wire  _T_30 = _T_29 | realDirty_23; // @[DataCache.scala 69:37]
  wire  _T_31 = _T_30 | realDirty_24; // @[DataCache.scala 69:37]
  wire  _T_32 = _T_31 | realDirty_25; // @[DataCache.scala 69:37]
  wire  _T_33 = _T_32 | realDirty_26; // @[DataCache.scala 69:37]
  wire  _T_34 = _T_33 | realDirty_27; // @[DataCache.scala 69:37]
  wire  _T_35 = _T_34 | realDirty_28; // @[DataCache.scala 69:37]
  wire  _T_36 = _T_35 | realDirty_29; // @[DataCache.scala 69:37]
  wire  _T_37 = _T_36 | realDirty_30; // @[DataCache.scala 69:37]
  wire  _T_38 = _T_37 | realDirty_31; // @[DataCache.scala 69:37]
  wire  _T_39 = _T_38 | realDirty_32; // @[DataCache.scala 69:37]
  wire  _T_40 = _T_39 | realDirty_33; // @[DataCache.scala 69:37]
  wire  _T_41 = _T_40 | realDirty_34; // @[DataCache.scala 69:37]
  wire  _T_42 = _T_41 | realDirty_35; // @[DataCache.scala 69:37]
  wire  _T_43 = _T_42 | realDirty_36; // @[DataCache.scala 69:37]
  wire  _T_44 = _T_43 | realDirty_37; // @[DataCache.scala 69:37]
  wire  _T_45 = _T_44 | realDirty_38; // @[DataCache.scala 69:37]
  wire  _T_46 = _T_45 | realDirty_39; // @[DataCache.scala 69:37]
  wire  _T_47 = _T_46 | realDirty_40; // @[DataCache.scala 69:37]
  wire  _T_48 = _T_47 | realDirty_41; // @[DataCache.scala 69:37]
  wire  _T_49 = _T_48 | realDirty_42; // @[DataCache.scala 69:37]
  wire  _T_50 = _T_49 | realDirty_43; // @[DataCache.scala 69:37]
  wire  _T_51 = _T_50 | realDirty_44; // @[DataCache.scala 69:37]
  wire  _T_52 = _T_51 | realDirty_45; // @[DataCache.scala 69:37]
  wire  _T_53 = _T_52 | realDirty_46; // @[DataCache.scala 69:37]
  wire  _T_54 = _T_53 | realDirty_47; // @[DataCache.scala 69:37]
  wire  _T_55 = _T_54 | realDirty_48; // @[DataCache.scala 69:37]
  wire  _T_56 = _T_55 | realDirty_49; // @[DataCache.scala 69:37]
  wire  _T_57 = _T_56 | realDirty_50; // @[DataCache.scala 69:37]
  wire  _T_58 = _T_57 | realDirty_51; // @[DataCache.scala 69:37]
  wire  _T_59 = _T_58 | realDirty_52; // @[DataCache.scala 69:37]
  wire  _T_60 = _T_59 | realDirty_53; // @[DataCache.scala 69:37]
  wire  _T_61 = _T_60 | realDirty_54; // @[DataCache.scala 69:37]
  wire  _T_62 = _T_61 | realDirty_55; // @[DataCache.scala 69:37]
  wire  _T_63 = _T_62 | realDirty_56; // @[DataCache.scala 69:37]
  wire  _T_64 = _T_63 | realDirty_57; // @[DataCache.scala 69:37]
  wire  _T_65 = _T_64 | realDirty_58; // @[DataCache.scala 69:37]
  wire  _T_66 = _T_65 | realDirty_59; // @[DataCache.scala 69:37]
  wire  _T_67 = _T_66 | realDirty_60; // @[DataCache.scala 69:37]
  wire  _T_68 = _T_67 | realDirty_61; // @[DataCache.scala 69:37]
  wire  _T_69 = _T_68 | realDirty_62; // @[DataCache.scala 69:37]
  wire  _T_70 = _T_69 | realDirty_63; // @[DataCache.scala 69:37]
  wire  _T_71 = _T_70 | realDirty_64; // @[DataCache.scala 69:37]
  wire  _T_72 = _T_71 | realDirty_65; // @[DataCache.scala 69:37]
  wire  _T_73 = _T_72 | realDirty_66; // @[DataCache.scala 69:37]
  wire  _T_74 = _T_73 | realDirty_67; // @[DataCache.scala 69:37]
  wire  _T_75 = _T_74 | realDirty_68; // @[DataCache.scala 69:37]
  wire  _T_76 = _T_75 | realDirty_69; // @[DataCache.scala 69:37]
  wire  _T_77 = _T_76 | realDirty_70; // @[DataCache.scala 69:37]
  wire  _T_78 = _T_77 | realDirty_71; // @[DataCache.scala 69:37]
  wire  _T_79 = _T_78 | realDirty_72; // @[DataCache.scala 69:37]
  wire  _T_80 = _T_79 | realDirty_73; // @[DataCache.scala 69:37]
  wire  _T_81 = _T_80 | realDirty_74; // @[DataCache.scala 69:37]
  wire  _T_82 = _T_81 | realDirty_75; // @[DataCache.scala 69:37]
  wire  _T_83 = _T_82 | realDirty_76; // @[DataCache.scala 69:37]
  wire  _T_84 = _T_83 | realDirty_77; // @[DataCache.scala 69:37]
  wire  _T_85 = _T_84 | realDirty_78; // @[DataCache.scala 69:37]
  wire  _T_86 = _T_85 | realDirty_79; // @[DataCache.scala 69:37]
  wire  _T_87 = _T_86 | realDirty_80; // @[DataCache.scala 69:37]
  wire  _T_88 = _T_87 | realDirty_81; // @[DataCache.scala 69:37]
  wire  _T_89 = _T_88 | realDirty_82; // @[DataCache.scala 69:37]
  wire  _T_90 = _T_89 | realDirty_83; // @[DataCache.scala 69:37]
  wire  _T_91 = _T_90 | realDirty_84; // @[DataCache.scala 69:37]
  wire  _T_92 = _T_91 | realDirty_85; // @[DataCache.scala 69:37]
  wire  _T_93 = _T_92 | realDirty_86; // @[DataCache.scala 69:37]
  wire  _T_94 = _T_93 | realDirty_87; // @[DataCache.scala 69:37]
  wire  _T_95 = _T_94 | realDirty_88; // @[DataCache.scala 69:37]
  wire  _T_96 = _T_95 | realDirty_89; // @[DataCache.scala 69:37]
  wire  _T_97 = _T_96 | realDirty_90; // @[DataCache.scala 69:37]
  wire  _T_98 = _T_97 | realDirty_91; // @[DataCache.scala 69:37]
  wire  _T_99 = _T_98 | realDirty_92; // @[DataCache.scala 69:37]
  wire  _T_100 = _T_99 | realDirty_93; // @[DataCache.scala 69:37]
  wire  _T_101 = _T_100 | realDirty_94; // @[DataCache.scala 69:37]
  wire  _T_102 = _T_101 | realDirty_95; // @[DataCache.scala 69:37]
  wire  _T_103 = _T_102 | realDirty_96; // @[DataCache.scala 69:37]
  wire  _T_104 = _T_103 | realDirty_97; // @[DataCache.scala 69:37]
  wire  _T_105 = _T_104 | realDirty_98; // @[DataCache.scala 69:37]
  wire  _T_106 = _T_105 | realDirty_99; // @[DataCache.scala 69:37]
  wire  _T_107 = _T_106 | realDirty_100; // @[DataCache.scala 69:37]
  wire  _T_108 = _T_107 | realDirty_101; // @[DataCache.scala 69:37]
  wire  _T_109 = _T_108 | realDirty_102; // @[DataCache.scala 69:37]
  wire  _T_110 = _T_109 | realDirty_103; // @[DataCache.scala 69:37]
  wire  _T_111 = _T_110 | realDirty_104; // @[DataCache.scala 69:37]
  wire  _T_112 = _T_111 | realDirty_105; // @[DataCache.scala 69:37]
  wire  _T_113 = _T_112 | realDirty_106; // @[DataCache.scala 69:37]
  wire  _T_114 = _T_113 | realDirty_107; // @[DataCache.scala 69:37]
  wire  _T_115 = _T_114 | realDirty_108; // @[DataCache.scala 69:37]
  wire  _T_116 = _T_115 | realDirty_109; // @[DataCache.scala 69:37]
  wire  _T_117 = _T_116 | realDirty_110; // @[DataCache.scala 69:37]
  wire  _T_118 = _T_117 | realDirty_111; // @[DataCache.scala 69:37]
  wire  _T_119 = _T_118 | realDirty_112; // @[DataCache.scala 69:37]
  wire  _T_120 = _T_119 | realDirty_113; // @[DataCache.scala 69:37]
  wire  _T_121 = _T_120 | realDirty_114; // @[DataCache.scala 69:37]
  wire  _T_122 = _T_121 | realDirty_115; // @[DataCache.scala 69:37]
  wire  _T_123 = _T_122 | realDirty_116; // @[DataCache.scala 69:37]
  wire  _T_124 = _T_123 | realDirty_117; // @[DataCache.scala 69:37]
  wire  _T_125 = _T_124 | realDirty_118; // @[DataCache.scala 69:37]
  wire  _T_126 = _T_125 | realDirty_119; // @[DataCache.scala 69:37]
  wire  _T_127 = _T_126 | realDirty_120; // @[DataCache.scala 69:37]
  wire  _T_128 = _T_127 | realDirty_121; // @[DataCache.scala 69:37]
  wire  _T_129 = _T_128 | realDirty_122; // @[DataCache.scala 69:37]
  wire  _T_130 = _T_129 | realDirty_123; // @[DataCache.scala 69:37]
  wire  _T_131 = _T_130 | realDirty_124; // @[DataCache.scala 69:37]
  wire  _T_132 = _T_131 | realDirty_125; // @[DataCache.scala 69:37]
  wire  _T_133 = _T_132 | realDirty_126; // @[DataCache.scala 69:37]
  wire  isDirty = _T_133 | realDirty_127; // @[DataCache.scala 69:37]
  wire [6:0] _T_134 = realDirty_126 ? 7'h7e : 7'h7f; // @[Mux.scala 47:69]
  wire [6:0] _T_135 = realDirty_125 ? 7'h7d : _T_134; // @[Mux.scala 47:69]
  wire [6:0] _T_136 = realDirty_124 ? 7'h7c : _T_135; // @[Mux.scala 47:69]
  wire [6:0] _T_137 = realDirty_123 ? 7'h7b : _T_136; // @[Mux.scala 47:69]
  wire [6:0] _T_138 = realDirty_122 ? 7'h7a : _T_137; // @[Mux.scala 47:69]
  wire [6:0] _T_139 = realDirty_121 ? 7'h79 : _T_138; // @[Mux.scala 47:69]
  wire [6:0] _T_140 = realDirty_120 ? 7'h78 : _T_139; // @[Mux.scala 47:69]
  wire [6:0] _T_141 = realDirty_119 ? 7'h77 : _T_140; // @[Mux.scala 47:69]
  wire [6:0] _T_142 = realDirty_118 ? 7'h76 : _T_141; // @[Mux.scala 47:69]
  wire [6:0] _T_143 = realDirty_117 ? 7'h75 : _T_142; // @[Mux.scala 47:69]
  wire [6:0] _T_144 = realDirty_116 ? 7'h74 : _T_143; // @[Mux.scala 47:69]
  wire [6:0] _T_145 = realDirty_115 ? 7'h73 : _T_144; // @[Mux.scala 47:69]
  wire [6:0] _T_146 = realDirty_114 ? 7'h72 : _T_145; // @[Mux.scala 47:69]
  wire [6:0] _T_147 = realDirty_113 ? 7'h71 : _T_146; // @[Mux.scala 47:69]
  wire [6:0] _T_148 = realDirty_112 ? 7'h70 : _T_147; // @[Mux.scala 47:69]
  wire [6:0] _T_149 = realDirty_111 ? 7'h6f : _T_148; // @[Mux.scala 47:69]
  wire [6:0] _T_150 = realDirty_110 ? 7'h6e : _T_149; // @[Mux.scala 47:69]
  wire [6:0] _T_151 = realDirty_109 ? 7'h6d : _T_150; // @[Mux.scala 47:69]
  wire [6:0] _T_152 = realDirty_108 ? 7'h6c : _T_151; // @[Mux.scala 47:69]
  wire [6:0] _T_153 = realDirty_107 ? 7'h6b : _T_152; // @[Mux.scala 47:69]
  wire [6:0] _T_154 = realDirty_106 ? 7'h6a : _T_153; // @[Mux.scala 47:69]
  wire [6:0] _T_155 = realDirty_105 ? 7'h69 : _T_154; // @[Mux.scala 47:69]
  wire [6:0] _T_156 = realDirty_104 ? 7'h68 : _T_155; // @[Mux.scala 47:69]
  wire [6:0] _T_157 = realDirty_103 ? 7'h67 : _T_156; // @[Mux.scala 47:69]
  wire [6:0] _T_158 = realDirty_102 ? 7'h66 : _T_157; // @[Mux.scala 47:69]
  wire [6:0] _T_159 = realDirty_101 ? 7'h65 : _T_158; // @[Mux.scala 47:69]
  wire [6:0] _T_160 = realDirty_100 ? 7'h64 : _T_159; // @[Mux.scala 47:69]
  wire [6:0] _T_161 = realDirty_99 ? 7'h63 : _T_160; // @[Mux.scala 47:69]
  wire [6:0] _T_162 = realDirty_98 ? 7'h62 : _T_161; // @[Mux.scala 47:69]
  wire [6:0] _T_163 = realDirty_97 ? 7'h61 : _T_162; // @[Mux.scala 47:69]
  wire [6:0] _T_164 = realDirty_96 ? 7'h60 : _T_163; // @[Mux.scala 47:69]
  wire [6:0] _T_165 = realDirty_95 ? 7'h5f : _T_164; // @[Mux.scala 47:69]
  wire [6:0] _T_166 = realDirty_94 ? 7'h5e : _T_165; // @[Mux.scala 47:69]
  wire [6:0] _T_167 = realDirty_93 ? 7'h5d : _T_166; // @[Mux.scala 47:69]
  wire [6:0] _T_168 = realDirty_92 ? 7'h5c : _T_167; // @[Mux.scala 47:69]
  wire [6:0] _T_169 = realDirty_91 ? 7'h5b : _T_168; // @[Mux.scala 47:69]
  wire [6:0] _T_170 = realDirty_90 ? 7'h5a : _T_169; // @[Mux.scala 47:69]
  wire [6:0] _T_171 = realDirty_89 ? 7'h59 : _T_170; // @[Mux.scala 47:69]
  wire [6:0] _T_172 = realDirty_88 ? 7'h58 : _T_171; // @[Mux.scala 47:69]
  wire [6:0] _T_173 = realDirty_87 ? 7'h57 : _T_172; // @[Mux.scala 47:69]
  wire [6:0] _T_174 = realDirty_86 ? 7'h56 : _T_173; // @[Mux.scala 47:69]
  wire [6:0] _T_175 = realDirty_85 ? 7'h55 : _T_174; // @[Mux.scala 47:69]
  wire [6:0] _T_176 = realDirty_84 ? 7'h54 : _T_175; // @[Mux.scala 47:69]
  wire [6:0] _T_177 = realDirty_83 ? 7'h53 : _T_176; // @[Mux.scala 47:69]
  wire [6:0] _T_178 = realDirty_82 ? 7'h52 : _T_177; // @[Mux.scala 47:69]
  wire [6:0] _T_179 = realDirty_81 ? 7'h51 : _T_178; // @[Mux.scala 47:69]
  wire [6:0] _T_180 = realDirty_80 ? 7'h50 : _T_179; // @[Mux.scala 47:69]
  wire [6:0] _T_181 = realDirty_79 ? 7'h4f : _T_180; // @[Mux.scala 47:69]
  wire [6:0] _T_182 = realDirty_78 ? 7'h4e : _T_181; // @[Mux.scala 47:69]
  wire [6:0] _T_183 = realDirty_77 ? 7'h4d : _T_182; // @[Mux.scala 47:69]
  wire [6:0] _T_184 = realDirty_76 ? 7'h4c : _T_183; // @[Mux.scala 47:69]
  wire [6:0] _T_185 = realDirty_75 ? 7'h4b : _T_184; // @[Mux.scala 47:69]
  wire [6:0] _T_186 = realDirty_74 ? 7'h4a : _T_185; // @[Mux.scala 47:69]
  wire [6:0] _T_187 = realDirty_73 ? 7'h49 : _T_186; // @[Mux.scala 47:69]
  wire [6:0] _T_188 = realDirty_72 ? 7'h48 : _T_187; // @[Mux.scala 47:69]
  wire [6:0] _T_189 = realDirty_71 ? 7'h47 : _T_188; // @[Mux.scala 47:69]
  wire [6:0] _T_190 = realDirty_70 ? 7'h46 : _T_189; // @[Mux.scala 47:69]
  wire [6:0] _T_191 = realDirty_69 ? 7'h45 : _T_190; // @[Mux.scala 47:69]
  wire [6:0] _T_192 = realDirty_68 ? 7'h44 : _T_191; // @[Mux.scala 47:69]
  wire [6:0] _T_193 = realDirty_67 ? 7'h43 : _T_192; // @[Mux.scala 47:69]
  wire [6:0] _T_194 = realDirty_66 ? 7'h42 : _T_193; // @[Mux.scala 47:69]
  wire [6:0] _T_195 = realDirty_65 ? 7'h41 : _T_194; // @[Mux.scala 47:69]
  wire [6:0] _T_196 = realDirty_64 ? 7'h40 : _T_195; // @[Mux.scala 47:69]
  wire [6:0] _T_197 = realDirty_63 ? 7'h3f : _T_196; // @[Mux.scala 47:69]
  wire [6:0] _T_198 = realDirty_62 ? 7'h3e : _T_197; // @[Mux.scala 47:69]
  wire [6:0] _T_199 = realDirty_61 ? 7'h3d : _T_198; // @[Mux.scala 47:69]
  wire [6:0] _T_200 = realDirty_60 ? 7'h3c : _T_199; // @[Mux.scala 47:69]
  wire [6:0] _T_201 = realDirty_59 ? 7'h3b : _T_200; // @[Mux.scala 47:69]
  wire [6:0] _T_202 = realDirty_58 ? 7'h3a : _T_201; // @[Mux.scala 47:69]
  wire [6:0] _T_203 = realDirty_57 ? 7'h39 : _T_202; // @[Mux.scala 47:69]
  wire [6:0] _T_204 = realDirty_56 ? 7'h38 : _T_203; // @[Mux.scala 47:69]
  wire [6:0] _T_205 = realDirty_55 ? 7'h37 : _T_204; // @[Mux.scala 47:69]
  wire [6:0] _T_206 = realDirty_54 ? 7'h36 : _T_205; // @[Mux.scala 47:69]
  wire [6:0] _T_207 = realDirty_53 ? 7'h35 : _T_206; // @[Mux.scala 47:69]
  wire [6:0] _T_208 = realDirty_52 ? 7'h34 : _T_207; // @[Mux.scala 47:69]
  wire [6:0] _T_209 = realDirty_51 ? 7'h33 : _T_208; // @[Mux.scala 47:69]
  wire [6:0] _T_210 = realDirty_50 ? 7'h32 : _T_209; // @[Mux.scala 47:69]
  wire [6:0] _T_211 = realDirty_49 ? 7'h31 : _T_210; // @[Mux.scala 47:69]
  wire [6:0] _T_212 = realDirty_48 ? 7'h30 : _T_211; // @[Mux.scala 47:69]
  wire [6:0] _T_213 = realDirty_47 ? 7'h2f : _T_212; // @[Mux.scala 47:69]
  wire [6:0] _T_214 = realDirty_46 ? 7'h2e : _T_213; // @[Mux.scala 47:69]
  wire [6:0] _T_215 = realDirty_45 ? 7'h2d : _T_214; // @[Mux.scala 47:69]
  wire [6:0] _T_216 = realDirty_44 ? 7'h2c : _T_215; // @[Mux.scala 47:69]
  wire [6:0] _T_217 = realDirty_43 ? 7'h2b : _T_216; // @[Mux.scala 47:69]
  wire [6:0] _T_218 = realDirty_42 ? 7'h2a : _T_217; // @[Mux.scala 47:69]
  wire [6:0] _T_219 = realDirty_41 ? 7'h29 : _T_218; // @[Mux.scala 47:69]
  wire [6:0] _T_220 = realDirty_40 ? 7'h28 : _T_219; // @[Mux.scala 47:69]
  wire [6:0] _T_221 = realDirty_39 ? 7'h27 : _T_220; // @[Mux.scala 47:69]
  wire [6:0] _T_222 = realDirty_38 ? 7'h26 : _T_221; // @[Mux.scala 47:69]
  wire [6:0] _T_223 = realDirty_37 ? 7'h25 : _T_222; // @[Mux.scala 47:69]
  wire [6:0] _T_224 = realDirty_36 ? 7'h24 : _T_223; // @[Mux.scala 47:69]
  wire [6:0] _T_225 = realDirty_35 ? 7'h23 : _T_224; // @[Mux.scala 47:69]
  wire [6:0] _T_226 = realDirty_34 ? 7'h22 : _T_225; // @[Mux.scala 47:69]
  wire [6:0] _T_227 = realDirty_33 ? 7'h21 : _T_226; // @[Mux.scala 47:69]
  wire [6:0] _T_228 = realDirty_32 ? 7'h20 : _T_227; // @[Mux.scala 47:69]
  wire [6:0] _T_229 = realDirty_31 ? 7'h1f : _T_228; // @[Mux.scala 47:69]
  wire [6:0] _T_230 = realDirty_30 ? 7'h1e : _T_229; // @[Mux.scala 47:69]
  wire [6:0] _T_231 = realDirty_29 ? 7'h1d : _T_230; // @[Mux.scala 47:69]
  wire [6:0] _T_232 = realDirty_28 ? 7'h1c : _T_231; // @[Mux.scala 47:69]
  wire [6:0] _T_233 = realDirty_27 ? 7'h1b : _T_232; // @[Mux.scala 47:69]
  wire [6:0] _T_234 = realDirty_26 ? 7'h1a : _T_233; // @[Mux.scala 47:69]
  wire [6:0] _T_235 = realDirty_25 ? 7'h19 : _T_234; // @[Mux.scala 47:69]
  wire [6:0] _T_236 = realDirty_24 ? 7'h18 : _T_235; // @[Mux.scala 47:69]
  wire [6:0] _T_237 = realDirty_23 ? 7'h17 : _T_236; // @[Mux.scala 47:69]
  wire [6:0] _T_238 = realDirty_22 ? 7'h16 : _T_237; // @[Mux.scala 47:69]
  wire [6:0] _T_239 = realDirty_21 ? 7'h15 : _T_238; // @[Mux.scala 47:69]
  wire [6:0] _T_240 = realDirty_20 ? 7'h14 : _T_239; // @[Mux.scala 47:69]
  wire [6:0] _T_241 = realDirty_19 ? 7'h13 : _T_240; // @[Mux.scala 47:69]
  wire [6:0] _T_242 = realDirty_18 ? 7'h12 : _T_241; // @[Mux.scala 47:69]
  wire [6:0] _T_243 = realDirty_17 ? 7'h11 : _T_242; // @[Mux.scala 47:69]
  wire [6:0] _T_244 = realDirty_16 ? 7'h10 : _T_243; // @[Mux.scala 47:69]
  wire [6:0] _T_245 = realDirty_15 ? 7'hf : _T_244; // @[Mux.scala 47:69]
  wire [6:0] _T_246 = realDirty_14 ? 7'he : _T_245; // @[Mux.scala 47:69]
  wire [6:0] _T_247 = realDirty_13 ? 7'hd : _T_246; // @[Mux.scala 47:69]
  wire [6:0] _T_248 = realDirty_12 ? 7'hc : _T_247; // @[Mux.scala 47:69]
  wire [6:0] _T_249 = realDirty_11 ? 7'hb : _T_248; // @[Mux.scala 47:69]
  wire [6:0] _T_250 = realDirty_10 ? 7'ha : _T_249; // @[Mux.scala 47:69]
  wire [6:0] _T_251 = realDirty_9 ? 7'h9 : _T_250; // @[Mux.scala 47:69]
  wire [6:0] _T_252 = realDirty_8 ? 7'h8 : _T_251; // @[Mux.scala 47:69]
  wire [6:0] _T_253 = realDirty_7 ? 7'h7 : _T_252; // @[Mux.scala 47:69]
  wire [6:0] _T_254 = realDirty_6 ? 7'h6 : _T_253; // @[Mux.scala 47:69]
  wire [6:0] _T_255 = realDirty_5 ? 7'h5 : _T_254; // @[Mux.scala 47:69]
  wire [6:0] _T_256 = realDirty_4 ? 7'h4 : _T_255; // @[Mux.scala 47:69]
  wire [6:0] _T_257 = realDirty_3 ? 7'h3 : _T_256; // @[Mux.scala 47:69]
  wire [6:0] _T_258 = realDirty_2 ? 7'h2 : _T_257; // @[Mux.scala 47:69]
  wire [6:0] _T_259 = realDirty_1 ? 7'h1 : _T_258; // @[Mux.scala 47:69]
  wire [6:0] nextDirty = realDirty_0 ? 7'h0 : _T_259; // @[Mux.scala 47:69]
  wire [31:0] flushAddr = {tag__T_261_data,nextDirty,6'h0}; // @[Cat.scala 30:58]
  wire [10:0] flushSel = {nextDirty,dataOfsRef}; // @[Cat.scala 30:58]
  wire  _T_264 = ~io_flush; // @[DataCache.scala 75:40]
  wire  _T_265 = _T_2 & _T_264; // @[DataCache.scala 75:37]
  wire  _T_266 = _T_265 & io_sram_en; // @[DataCache.scala 75:50]
  wire  lineEnCpu = _T_266 & cacheHit; // @[DataCache.scala 75:64]
  wire  _T_267 = state == 4'h2; // @[DataCache.scala 76:27]
  wire  lineEnRead = _T_267 & io_axi_readData_valid; // @[DataCache.scala 76:41]
  wire  lineEnWrite = state == 4'h5; // @[DataCache.scala 77:27]
  wire  lineEnFlush = state == 4'h7; // @[DataCache.scala 78:27]
  wire [3:0] _T_268 = lineEnRead ? 4'hf : 4'h0; // @[DataCache.scala 81:25]
  wire  _T_270 = lineEnRead | lineEnWrite; // @[DataCache.scala 82:37]
  wire [10:0] _T_271 = lineEnFlush ? flushSel : lineDataSel; // @[DataCache.scala 83:25]
  wire  _T_274 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_275 = io_flush & isDirty; // @[DataCache.scala 91:22]
  wire  _T_276 = io_sram_wen != 4'h0; // @[DataCache.scala 97:29]
  wire  _GEN_3427 = 7'h0 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_128 = _GEN_3427 | dirty_0; // @[DataCache.scala 99:28]
  wire  _GEN_3428 = 7'h1 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_129 = _GEN_3428 | dirty_1; // @[DataCache.scala 99:28]
  wire  _GEN_3429 = 7'h2 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_130 = _GEN_3429 | dirty_2; // @[DataCache.scala 99:28]
  wire  _GEN_3430 = 7'h3 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_131 = _GEN_3430 | dirty_3; // @[DataCache.scala 99:28]
  wire  _GEN_3431 = 7'h4 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_132 = _GEN_3431 | dirty_4; // @[DataCache.scala 99:28]
  wire  _GEN_3432 = 7'h5 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_133 = _GEN_3432 | dirty_5; // @[DataCache.scala 99:28]
  wire  _GEN_3433 = 7'h6 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_134 = _GEN_3433 | dirty_6; // @[DataCache.scala 99:28]
  wire  _GEN_3434 = 7'h7 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_135 = _GEN_3434 | dirty_7; // @[DataCache.scala 99:28]
  wire  _GEN_3435 = 7'h8 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_136 = _GEN_3435 | dirty_8; // @[DataCache.scala 99:28]
  wire  _GEN_3436 = 7'h9 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_137 = _GEN_3436 | dirty_9; // @[DataCache.scala 99:28]
  wire  _GEN_3437 = 7'ha == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_138 = _GEN_3437 | dirty_10; // @[DataCache.scala 99:28]
  wire  _GEN_3438 = 7'hb == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_139 = _GEN_3438 | dirty_11; // @[DataCache.scala 99:28]
  wire  _GEN_3439 = 7'hc == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_140 = _GEN_3439 | dirty_12; // @[DataCache.scala 99:28]
  wire  _GEN_3440 = 7'hd == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_141 = _GEN_3440 | dirty_13; // @[DataCache.scala 99:28]
  wire  _GEN_3441 = 7'he == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_142 = _GEN_3441 | dirty_14; // @[DataCache.scala 99:28]
  wire  _GEN_3442 = 7'hf == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_143 = _GEN_3442 | dirty_15; // @[DataCache.scala 99:28]
  wire  _GEN_3443 = 7'h10 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_144 = _GEN_3443 | dirty_16; // @[DataCache.scala 99:28]
  wire  _GEN_3444 = 7'h11 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_145 = _GEN_3444 | dirty_17; // @[DataCache.scala 99:28]
  wire  _GEN_3445 = 7'h12 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_146 = _GEN_3445 | dirty_18; // @[DataCache.scala 99:28]
  wire  _GEN_3446 = 7'h13 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_147 = _GEN_3446 | dirty_19; // @[DataCache.scala 99:28]
  wire  _GEN_3447 = 7'h14 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_148 = _GEN_3447 | dirty_20; // @[DataCache.scala 99:28]
  wire  _GEN_3448 = 7'h15 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_149 = _GEN_3448 | dirty_21; // @[DataCache.scala 99:28]
  wire  _GEN_3449 = 7'h16 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_150 = _GEN_3449 | dirty_22; // @[DataCache.scala 99:28]
  wire  _GEN_3450 = 7'h17 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_151 = _GEN_3450 | dirty_23; // @[DataCache.scala 99:28]
  wire  _GEN_3451 = 7'h18 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_152 = _GEN_3451 | dirty_24; // @[DataCache.scala 99:28]
  wire  _GEN_3452 = 7'h19 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_153 = _GEN_3452 | dirty_25; // @[DataCache.scala 99:28]
  wire  _GEN_3453 = 7'h1a == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_154 = _GEN_3453 | dirty_26; // @[DataCache.scala 99:28]
  wire  _GEN_3454 = 7'h1b == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_155 = _GEN_3454 | dirty_27; // @[DataCache.scala 99:28]
  wire  _GEN_3455 = 7'h1c == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_156 = _GEN_3455 | dirty_28; // @[DataCache.scala 99:28]
  wire  _GEN_3456 = 7'h1d == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_157 = _GEN_3456 | dirty_29; // @[DataCache.scala 99:28]
  wire  _GEN_3457 = 7'h1e == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_158 = _GEN_3457 | dirty_30; // @[DataCache.scala 99:28]
  wire  _GEN_3458 = 7'h1f == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_159 = _GEN_3458 | dirty_31; // @[DataCache.scala 99:28]
  wire  _GEN_3459 = 7'h20 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_160 = _GEN_3459 | dirty_32; // @[DataCache.scala 99:28]
  wire  _GEN_3460 = 7'h21 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_161 = _GEN_3460 | dirty_33; // @[DataCache.scala 99:28]
  wire  _GEN_3461 = 7'h22 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_162 = _GEN_3461 | dirty_34; // @[DataCache.scala 99:28]
  wire  _GEN_3462 = 7'h23 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_163 = _GEN_3462 | dirty_35; // @[DataCache.scala 99:28]
  wire  _GEN_3463 = 7'h24 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_164 = _GEN_3463 | dirty_36; // @[DataCache.scala 99:28]
  wire  _GEN_3464 = 7'h25 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_165 = _GEN_3464 | dirty_37; // @[DataCache.scala 99:28]
  wire  _GEN_3465 = 7'h26 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_166 = _GEN_3465 | dirty_38; // @[DataCache.scala 99:28]
  wire  _GEN_3466 = 7'h27 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_167 = _GEN_3466 | dirty_39; // @[DataCache.scala 99:28]
  wire  _GEN_3467 = 7'h28 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_168 = _GEN_3467 | dirty_40; // @[DataCache.scala 99:28]
  wire  _GEN_3468 = 7'h29 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_169 = _GEN_3468 | dirty_41; // @[DataCache.scala 99:28]
  wire  _GEN_3469 = 7'h2a == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_170 = _GEN_3469 | dirty_42; // @[DataCache.scala 99:28]
  wire  _GEN_3470 = 7'h2b == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_171 = _GEN_3470 | dirty_43; // @[DataCache.scala 99:28]
  wire  _GEN_3471 = 7'h2c == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_172 = _GEN_3471 | dirty_44; // @[DataCache.scala 99:28]
  wire  _GEN_3472 = 7'h2d == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_173 = _GEN_3472 | dirty_45; // @[DataCache.scala 99:28]
  wire  _GEN_3473 = 7'h2e == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_174 = _GEN_3473 | dirty_46; // @[DataCache.scala 99:28]
  wire  _GEN_3474 = 7'h2f == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_175 = _GEN_3474 | dirty_47; // @[DataCache.scala 99:28]
  wire  _GEN_3475 = 7'h30 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_176 = _GEN_3475 | dirty_48; // @[DataCache.scala 99:28]
  wire  _GEN_3476 = 7'h31 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_177 = _GEN_3476 | dirty_49; // @[DataCache.scala 99:28]
  wire  _GEN_3477 = 7'h32 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_178 = _GEN_3477 | dirty_50; // @[DataCache.scala 99:28]
  wire  _GEN_3478 = 7'h33 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_179 = _GEN_3478 | dirty_51; // @[DataCache.scala 99:28]
  wire  _GEN_3479 = 7'h34 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_180 = _GEN_3479 | dirty_52; // @[DataCache.scala 99:28]
  wire  _GEN_3480 = 7'h35 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_181 = _GEN_3480 | dirty_53; // @[DataCache.scala 99:28]
  wire  _GEN_3481 = 7'h36 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_182 = _GEN_3481 | dirty_54; // @[DataCache.scala 99:28]
  wire  _GEN_3482 = 7'h37 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_183 = _GEN_3482 | dirty_55; // @[DataCache.scala 99:28]
  wire  _GEN_3483 = 7'h38 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_184 = _GEN_3483 | dirty_56; // @[DataCache.scala 99:28]
  wire  _GEN_3484 = 7'h39 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_185 = _GEN_3484 | dirty_57; // @[DataCache.scala 99:28]
  wire  _GEN_3485 = 7'h3a == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_186 = _GEN_3485 | dirty_58; // @[DataCache.scala 99:28]
  wire  _GEN_3486 = 7'h3b == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_187 = _GEN_3486 | dirty_59; // @[DataCache.scala 99:28]
  wire  _GEN_3487 = 7'h3c == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_188 = _GEN_3487 | dirty_60; // @[DataCache.scala 99:28]
  wire  _GEN_3488 = 7'h3d == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_189 = _GEN_3488 | dirty_61; // @[DataCache.scala 99:28]
  wire  _GEN_3489 = 7'h3e == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_190 = _GEN_3489 | dirty_62; // @[DataCache.scala 99:28]
  wire  _GEN_3490 = 7'h3f == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_191 = _GEN_3490 | dirty_63; // @[DataCache.scala 99:28]
  wire  _GEN_3491 = 7'h40 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_192 = _GEN_3491 | dirty_64; // @[DataCache.scala 99:28]
  wire  _GEN_3492 = 7'h41 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_193 = _GEN_3492 | dirty_65; // @[DataCache.scala 99:28]
  wire  _GEN_3493 = 7'h42 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_194 = _GEN_3493 | dirty_66; // @[DataCache.scala 99:28]
  wire  _GEN_3494 = 7'h43 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_195 = _GEN_3494 | dirty_67; // @[DataCache.scala 99:28]
  wire  _GEN_3495 = 7'h44 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_196 = _GEN_3495 | dirty_68; // @[DataCache.scala 99:28]
  wire  _GEN_3496 = 7'h45 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_197 = _GEN_3496 | dirty_69; // @[DataCache.scala 99:28]
  wire  _GEN_3497 = 7'h46 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_198 = _GEN_3497 | dirty_70; // @[DataCache.scala 99:28]
  wire  _GEN_3498 = 7'h47 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_199 = _GEN_3498 | dirty_71; // @[DataCache.scala 99:28]
  wire  _GEN_3499 = 7'h48 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_200 = _GEN_3499 | dirty_72; // @[DataCache.scala 99:28]
  wire  _GEN_3500 = 7'h49 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_201 = _GEN_3500 | dirty_73; // @[DataCache.scala 99:28]
  wire  _GEN_3501 = 7'h4a == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_202 = _GEN_3501 | dirty_74; // @[DataCache.scala 99:28]
  wire  _GEN_3502 = 7'h4b == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_203 = _GEN_3502 | dirty_75; // @[DataCache.scala 99:28]
  wire  _GEN_3503 = 7'h4c == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_204 = _GEN_3503 | dirty_76; // @[DataCache.scala 99:28]
  wire  _GEN_3504 = 7'h4d == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_205 = _GEN_3504 | dirty_77; // @[DataCache.scala 99:28]
  wire  _GEN_3505 = 7'h4e == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_206 = _GEN_3505 | dirty_78; // @[DataCache.scala 99:28]
  wire  _GEN_3506 = 7'h4f == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_207 = _GEN_3506 | dirty_79; // @[DataCache.scala 99:28]
  wire  _GEN_3507 = 7'h50 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_208 = _GEN_3507 | dirty_80; // @[DataCache.scala 99:28]
  wire  _GEN_3508 = 7'h51 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_209 = _GEN_3508 | dirty_81; // @[DataCache.scala 99:28]
  wire  _GEN_3509 = 7'h52 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_210 = _GEN_3509 | dirty_82; // @[DataCache.scala 99:28]
  wire  _GEN_3510 = 7'h53 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_211 = _GEN_3510 | dirty_83; // @[DataCache.scala 99:28]
  wire  _GEN_3511 = 7'h54 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_212 = _GEN_3511 | dirty_84; // @[DataCache.scala 99:28]
  wire  _GEN_3512 = 7'h55 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_213 = _GEN_3512 | dirty_85; // @[DataCache.scala 99:28]
  wire  _GEN_3513 = 7'h56 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_214 = _GEN_3513 | dirty_86; // @[DataCache.scala 99:28]
  wire  _GEN_3514 = 7'h57 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_215 = _GEN_3514 | dirty_87; // @[DataCache.scala 99:28]
  wire  _GEN_3515 = 7'h58 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_216 = _GEN_3515 | dirty_88; // @[DataCache.scala 99:28]
  wire  _GEN_3516 = 7'h59 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_217 = _GEN_3516 | dirty_89; // @[DataCache.scala 99:28]
  wire  _GEN_3517 = 7'h5a == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_218 = _GEN_3517 | dirty_90; // @[DataCache.scala 99:28]
  wire  _GEN_3518 = 7'h5b == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_219 = _GEN_3518 | dirty_91; // @[DataCache.scala 99:28]
  wire  _GEN_3519 = 7'h5c == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_220 = _GEN_3519 | dirty_92; // @[DataCache.scala 99:28]
  wire  _GEN_3520 = 7'h5d == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_221 = _GEN_3520 | dirty_93; // @[DataCache.scala 99:28]
  wire  _GEN_3521 = 7'h5e == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_222 = _GEN_3521 | dirty_94; // @[DataCache.scala 99:28]
  wire  _GEN_3522 = 7'h5f == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_223 = _GEN_3522 | dirty_95; // @[DataCache.scala 99:28]
  wire  _GEN_3523 = 7'h60 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_224 = _GEN_3523 | dirty_96; // @[DataCache.scala 99:28]
  wire  _GEN_3524 = 7'h61 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_225 = _GEN_3524 | dirty_97; // @[DataCache.scala 99:28]
  wire  _GEN_3525 = 7'h62 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_226 = _GEN_3525 | dirty_98; // @[DataCache.scala 99:28]
  wire  _GEN_3526 = 7'h63 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_227 = _GEN_3526 | dirty_99; // @[DataCache.scala 99:28]
  wire  _GEN_3527 = 7'h64 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_228 = _GEN_3527 | dirty_100; // @[DataCache.scala 99:28]
  wire  _GEN_3528 = 7'h65 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_229 = _GEN_3528 | dirty_101; // @[DataCache.scala 99:28]
  wire  _GEN_3529 = 7'h66 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_230 = _GEN_3529 | dirty_102; // @[DataCache.scala 99:28]
  wire  _GEN_3530 = 7'h67 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_231 = _GEN_3530 | dirty_103; // @[DataCache.scala 99:28]
  wire  _GEN_3531 = 7'h68 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_232 = _GEN_3531 | dirty_104; // @[DataCache.scala 99:28]
  wire  _GEN_3532 = 7'h69 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_233 = _GEN_3532 | dirty_105; // @[DataCache.scala 99:28]
  wire  _GEN_3533 = 7'h6a == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_234 = _GEN_3533 | dirty_106; // @[DataCache.scala 99:28]
  wire  _GEN_3534 = 7'h6b == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_235 = _GEN_3534 | dirty_107; // @[DataCache.scala 99:28]
  wire  _GEN_3535 = 7'h6c == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_236 = _GEN_3535 | dirty_108; // @[DataCache.scala 99:28]
  wire  _GEN_3536 = 7'h6d == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_237 = _GEN_3536 | dirty_109; // @[DataCache.scala 99:28]
  wire  _GEN_3537 = 7'h6e == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_238 = _GEN_3537 | dirty_110; // @[DataCache.scala 99:28]
  wire  _GEN_3538 = 7'h6f == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_239 = _GEN_3538 | dirty_111; // @[DataCache.scala 99:28]
  wire  _GEN_3539 = 7'h70 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_240 = _GEN_3539 | dirty_112; // @[DataCache.scala 99:28]
  wire  _GEN_3540 = 7'h71 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_241 = _GEN_3540 | dirty_113; // @[DataCache.scala 99:28]
  wire  _GEN_3541 = 7'h72 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_242 = _GEN_3541 | dirty_114; // @[DataCache.scala 99:28]
  wire  _GEN_3542 = 7'h73 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_243 = _GEN_3542 | dirty_115; // @[DataCache.scala 99:28]
  wire  _GEN_3543 = 7'h74 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_244 = _GEN_3543 | dirty_116; // @[DataCache.scala 99:28]
  wire  _GEN_3544 = 7'h75 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_245 = _GEN_3544 | dirty_117; // @[DataCache.scala 99:28]
  wire  _GEN_3545 = 7'h76 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_246 = _GEN_3545 | dirty_118; // @[DataCache.scala 99:28]
  wire  _GEN_3546 = 7'h77 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_247 = _GEN_3546 | dirty_119; // @[DataCache.scala 99:28]
  wire  _GEN_3547 = 7'h78 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_248 = _GEN_3547 | dirty_120; // @[DataCache.scala 99:28]
  wire  _GEN_3548 = 7'h79 == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_249 = _GEN_3548 | dirty_121; // @[DataCache.scala 99:28]
  wire  _GEN_3549 = 7'h7a == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_250 = _GEN_3549 | dirty_122; // @[DataCache.scala 99:28]
  wire  _GEN_3550 = 7'h7b == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_251 = _GEN_3550 | dirty_123; // @[DataCache.scala 99:28]
  wire  _GEN_3551 = 7'h7c == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_252 = _GEN_3551 | dirty_124; // @[DataCache.scala 99:28]
  wire  _GEN_3552 = 7'h7d == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_253 = _GEN_3552 | dirty_125; // @[DataCache.scala 99:28]
  wire  _GEN_3553 = 7'h7e == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_254 = _GEN_3553 | dirty_126; // @[DataCache.scala 99:28]
  wire  _GEN_3554 = 7'h7f == lineSel; // @[DataCache.scala 99:28]
  wire  _GEN_255 = _GEN_3554 | dirty_127; // @[DataCache.scala 99:28]
  wire  _GEN_385 = 7'h1 == lineSel ? dirty_1 : dirty_0; // @[DataCache.scala 101:37]
  wire  _GEN_386 = 7'h2 == lineSel ? dirty_2 : _GEN_385; // @[DataCache.scala 101:37]
  wire  _GEN_387 = 7'h3 == lineSel ? dirty_3 : _GEN_386; // @[DataCache.scala 101:37]
  wire  _GEN_388 = 7'h4 == lineSel ? dirty_4 : _GEN_387; // @[DataCache.scala 101:37]
  wire  _GEN_389 = 7'h5 == lineSel ? dirty_5 : _GEN_388; // @[DataCache.scala 101:37]
  wire  _GEN_390 = 7'h6 == lineSel ? dirty_6 : _GEN_389; // @[DataCache.scala 101:37]
  wire  _GEN_391 = 7'h7 == lineSel ? dirty_7 : _GEN_390; // @[DataCache.scala 101:37]
  wire  _GEN_392 = 7'h8 == lineSel ? dirty_8 : _GEN_391; // @[DataCache.scala 101:37]
  wire  _GEN_393 = 7'h9 == lineSel ? dirty_9 : _GEN_392; // @[DataCache.scala 101:37]
  wire  _GEN_394 = 7'ha == lineSel ? dirty_10 : _GEN_393; // @[DataCache.scala 101:37]
  wire  _GEN_395 = 7'hb == lineSel ? dirty_11 : _GEN_394; // @[DataCache.scala 101:37]
  wire  _GEN_396 = 7'hc == lineSel ? dirty_12 : _GEN_395; // @[DataCache.scala 101:37]
  wire  _GEN_397 = 7'hd == lineSel ? dirty_13 : _GEN_396; // @[DataCache.scala 101:37]
  wire  _GEN_398 = 7'he == lineSel ? dirty_14 : _GEN_397; // @[DataCache.scala 101:37]
  wire  _GEN_399 = 7'hf == lineSel ? dirty_15 : _GEN_398; // @[DataCache.scala 101:37]
  wire  _GEN_400 = 7'h10 == lineSel ? dirty_16 : _GEN_399; // @[DataCache.scala 101:37]
  wire  _GEN_401 = 7'h11 == lineSel ? dirty_17 : _GEN_400; // @[DataCache.scala 101:37]
  wire  _GEN_402 = 7'h12 == lineSel ? dirty_18 : _GEN_401; // @[DataCache.scala 101:37]
  wire  _GEN_403 = 7'h13 == lineSel ? dirty_19 : _GEN_402; // @[DataCache.scala 101:37]
  wire  _GEN_404 = 7'h14 == lineSel ? dirty_20 : _GEN_403; // @[DataCache.scala 101:37]
  wire  _GEN_405 = 7'h15 == lineSel ? dirty_21 : _GEN_404; // @[DataCache.scala 101:37]
  wire  _GEN_406 = 7'h16 == lineSel ? dirty_22 : _GEN_405; // @[DataCache.scala 101:37]
  wire  _GEN_407 = 7'h17 == lineSel ? dirty_23 : _GEN_406; // @[DataCache.scala 101:37]
  wire  _GEN_408 = 7'h18 == lineSel ? dirty_24 : _GEN_407; // @[DataCache.scala 101:37]
  wire  _GEN_409 = 7'h19 == lineSel ? dirty_25 : _GEN_408; // @[DataCache.scala 101:37]
  wire  _GEN_410 = 7'h1a == lineSel ? dirty_26 : _GEN_409; // @[DataCache.scala 101:37]
  wire  _GEN_411 = 7'h1b == lineSel ? dirty_27 : _GEN_410; // @[DataCache.scala 101:37]
  wire  _GEN_412 = 7'h1c == lineSel ? dirty_28 : _GEN_411; // @[DataCache.scala 101:37]
  wire  _GEN_413 = 7'h1d == lineSel ? dirty_29 : _GEN_412; // @[DataCache.scala 101:37]
  wire  _GEN_414 = 7'h1e == lineSel ? dirty_30 : _GEN_413; // @[DataCache.scala 101:37]
  wire  _GEN_415 = 7'h1f == lineSel ? dirty_31 : _GEN_414; // @[DataCache.scala 101:37]
  wire  _GEN_416 = 7'h20 == lineSel ? dirty_32 : _GEN_415; // @[DataCache.scala 101:37]
  wire  _GEN_417 = 7'h21 == lineSel ? dirty_33 : _GEN_416; // @[DataCache.scala 101:37]
  wire  _GEN_418 = 7'h22 == lineSel ? dirty_34 : _GEN_417; // @[DataCache.scala 101:37]
  wire  _GEN_419 = 7'h23 == lineSel ? dirty_35 : _GEN_418; // @[DataCache.scala 101:37]
  wire  _GEN_420 = 7'h24 == lineSel ? dirty_36 : _GEN_419; // @[DataCache.scala 101:37]
  wire  _GEN_421 = 7'h25 == lineSel ? dirty_37 : _GEN_420; // @[DataCache.scala 101:37]
  wire  _GEN_422 = 7'h26 == lineSel ? dirty_38 : _GEN_421; // @[DataCache.scala 101:37]
  wire  _GEN_423 = 7'h27 == lineSel ? dirty_39 : _GEN_422; // @[DataCache.scala 101:37]
  wire  _GEN_424 = 7'h28 == lineSel ? dirty_40 : _GEN_423; // @[DataCache.scala 101:37]
  wire  _GEN_425 = 7'h29 == lineSel ? dirty_41 : _GEN_424; // @[DataCache.scala 101:37]
  wire  _GEN_426 = 7'h2a == lineSel ? dirty_42 : _GEN_425; // @[DataCache.scala 101:37]
  wire  _GEN_427 = 7'h2b == lineSel ? dirty_43 : _GEN_426; // @[DataCache.scala 101:37]
  wire  _GEN_428 = 7'h2c == lineSel ? dirty_44 : _GEN_427; // @[DataCache.scala 101:37]
  wire  _GEN_429 = 7'h2d == lineSel ? dirty_45 : _GEN_428; // @[DataCache.scala 101:37]
  wire  _GEN_430 = 7'h2e == lineSel ? dirty_46 : _GEN_429; // @[DataCache.scala 101:37]
  wire  _GEN_431 = 7'h2f == lineSel ? dirty_47 : _GEN_430; // @[DataCache.scala 101:37]
  wire  _GEN_432 = 7'h30 == lineSel ? dirty_48 : _GEN_431; // @[DataCache.scala 101:37]
  wire  _GEN_433 = 7'h31 == lineSel ? dirty_49 : _GEN_432; // @[DataCache.scala 101:37]
  wire  _GEN_434 = 7'h32 == lineSel ? dirty_50 : _GEN_433; // @[DataCache.scala 101:37]
  wire  _GEN_435 = 7'h33 == lineSel ? dirty_51 : _GEN_434; // @[DataCache.scala 101:37]
  wire  _GEN_436 = 7'h34 == lineSel ? dirty_52 : _GEN_435; // @[DataCache.scala 101:37]
  wire  _GEN_437 = 7'h35 == lineSel ? dirty_53 : _GEN_436; // @[DataCache.scala 101:37]
  wire  _GEN_438 = 7'h36 == lineSel ? dirty_54 : _GEN_437; // @[DataCache.scala 101:37]
  wire  _GEN_439 = 7'h37 == lineSel ? dirty_55 : _GEN_438; // @[DataCache.scala 101:37]
  wire  _GEN_440 = 7'h38 == lineSel ? dirty_56 : _GEN_439; // @[DataCache.scala 101:37]
  wire  _GEN_441 = 7'h39 == lineSel ? dirty_57 : _GEN_440; // @[DataCache.scala 101:37]
  wire  _GEN_442 = 7'h3a == lineSel ? dirty_58 : _GEN_441; // @[DataCache.scala 101:37]
  wire  _GEN_443 = 7'h3b == lineSel ? dirty_59 : _GEN_442; // @[DataCache.scala 101:37]
  wire  _GEN_444 = 7'h3c == lineSel ? dirty_60 : _GEN_443; // @[DataCache.scala 101:37]
  wire  _GEN_445 = 7'h3d == lineSel ? dirty_61 : _GEN_444; // @[DataCache.scala 101:37]
  wire  _GEN_446 = 7'h3e == lineSel ? dirty_62 : _GEN_445; // @[DataCache.scala 101:37]
  wire  _GEN_447 = 7'h3f == lineSel ? dirty_63 : _GEN_446; // @[DataCache.scala 101:37]
  wire  _GEN_448 = 7'h40 == lineSel ? dirty_64 : _GEN_447; // @[DataCache.scala 101:37]
  wire  _GEN_449 = 7'h41 == lineSel ? dirty_65 : _GEN_448; // @[DataCache.scala 101:37]
  wire  _GEN_450 = 7'h42 == lineSel ? dirty_66 : _GEN_449; // @[DataCache.scala 101:37]
  wire  _GEN_451 = 7'h43 == lineSel ? dirty_67 : _GEN_450; // @[DataCache.scala 101:37]
  wire  _GEN_452 = 7'h44 == lineSel ? dirty_68 : _GEN_451; // @[DataCache.scala 101:37]
  wire  _GEN_453 = 7'h45 == lineSel ? dirty_69 : _GEN_452; // @[DataCache.scala 101:37]
  wire  _GEN_454 = 7'h46 == lineSel ? dirty_70 : _GEN_453; // @[DataCache.scala 101:37]
  wire  _GEN_455 = 7'h47 == lineSel ? dirty_71 : _GEN_454; // @[DataCache.scala 101:37]
  wire  _GEN_456 = 7'h48 == lineSel ? dirty_72 : _GEN_455; // @[DataCache.scala 101:37]
  wire  _GEN_457 = 7'h49 == lineSel ? dirty_73 : _GEN_456; // @[DataCache.scala 101:37]
  wire  _GEN_458 = 7'h4a == lineSel ? dirty_74 : _GEN_457; // @[DataCache.scala 101:37]
  wire  _GEN_459 = 7'h4b == lineSel ? dirty_75 : _GEN_458; // @[DataCache.scala 101:37]
  wire  _GEN_460 = 7'h4c == lineSel ? dirty_76 : _GEN_459; // @[DataCache.scala 101:37]
  wire  _GEN_461 = 7'h4d == lineSel ? dirty_77 : _GEN_460; // @[DataCache.scala 101:37]
  wire  _GEN_462 = 7'h4e == lineSel ? dirty_78 : _GEN_461; // @[DataCache.scala 101:37]
  wire  _GEN_463 = 7'h4f == lineSel ? dirty_79 : _GEN_462; // @[DataCache.scala 101:37]
  wire  _GEN_464 = 7'h50 == lineSel ? dirty_80 : _GEN_463; // @[DataCache.scala 101:37]
  wire  _GEN_465 = 7'h51 == lineSel ? dirty_81 : _GEN_464; // @[DataCache.scala 101:37]
  wire  _GEN_466 = 7'h52 == lineSel ? dirty_82 : _GEN_465; // @[DataCache.scala 101:37]
  wire  _GEN_467 = 7'h53 == lineSel ? dirty_83 : _GEN_466; // @[DataCache.scala 101:37]
  wire  _GEN_468 = 7'h54 == lineSel ? dirty_84 : _GEN_467; // @[DataCache.scala 101:37]
  wire  _GEN_469 = 7'h55 == lineSel ? dirty_85 : _GEN_468; // @[DataCache.scala 101:37]
  wire  _GEN_470 = 7'h56 == lineSel ? dirty_86 : _GEN_469; // @[DataCache.scala 101:37]
  wire  _GEN_471 = 7'h57 == lineSel ? dirty_87 : _GEN_470; // @[DataCache.scala 101:37]
  wire  _GEN_472 = 7'h58 == lineSel ? dirty_88 : _GEN_471; // @[DataCache.scala 101:37]
  wire  _GEN_473 = 7'h59 == lineSel ? dirty_89 : _GEN_472; // @[DataCache.scala 101:37]
  wire  _GEN_474 = 7'h5a == lineSel ? dirty_90 : _GEN_473; // @[DataCache.scala 101:37]
  wire  _GEN_475 = 7'h5b == lineSel ? dirty_91 : _GEN_474; // @[DataCache.scala 101:37]
  wire  _GEN_476 = 7'h5c == lineSel ? dirty_92 : _GEN_475; // @[DataCache.scala 101:37]
  wire  _GEN_477 = 7'h5d == lineSel ? dirty_93 : _GEN_476; // @[DataCache.scala 101:37]
  wire  _GEN_478 = 7'h5e == lineSel ? dirty_94 : _GEN_477; // @[DataCache.scala 101:37]
  wire  _GEN_479 = 7'h5f == lineSel ? dirty_95 : _GEN_478; // @[DataCache.scala 101:37]
  wire  _GEN_480 = 7'h60 == lineSel ? dirty_96 : _GEN_479; // @[DataCache.scala 101:37]
  wire  _GEN_481 = 7'h61 == lineSel ? dirty_97 : _GEN_480; // @[DataCache.scala 101:37]
  wire  _GEN_482 = 7'h62 == lineSel ? dirty_98 : _GEN_481; // @[DataCache.scala 101:37]
  wire  _GEN_483 = 7'h63 == lineSel ? dirty_99 : _GEN_482; // @[DataCache.scala 101:37]
  wire  _GEN_484 = 7'h64 == lineSel ? dirty_100 : _GEN_483; // @[DataCache.scala 101:37]
  wire  _GEN_485 = 7'h65 == lineSel ? dirty_101 : _GEN_484; // @[DataCache.scala 101:37]
  wire  _GEN_486 = 7'h66 == lineSel ? dirty_102 : _GEN_485; // @[DataCache.scala 101:37]
  wire  _GEN_487 = 7'h67 == lineSel ? dirty_103 : _GEN_486; // @[DataCache.scala 101:37]
  wire  _GEN_488 = 7'h68 == lineSel ? dirty_104 : _GEN_487; // @[DataCache.scala 101:37]
  wire  _GEN_489 = 7'h69 == lineSel ? dirty_105 : _GEN_488; // @[DataCache.scala 101:37]
  wire  _GEN_490 = 7'h6a == lineSel ? dirty_106 : _GEN_489; // @[DataCache.scala 101:37]
  wire  _GEN_491 = 7'h6b == lineSel ? dirty_107 : _GEN_490; // @[DataCache.scala 101:37]
  wire  _GEN_492 = 7'h6c == lineSel ? dirty_108 : _GEN_491; // @[DataCache.scala 101:37]
  wire  _GEN_493 = 7'h6d == lineSel ? dirty_109 : _GEN_492; // @[DataCache.scala 101:37]
  wire  _GEN_494 = 7'h6e == lineSel ? dirty_110 : _GEN_493; // @[DataCache.scala 101:37]
  wire  _GEN_495 = 7'h6f == lineSel ? dirty_111 : _GEN_494; // @[DataCache.scala 101:37]
  wire  _GEN_496 = 7'h70 == lineSel ? dirty_112 : _GEN_495; // @[DataCache.scala 101:37]
  wire  _GEN_497 = 7'h71 == lineSel ? dirty_113 : _GEN_496; // @[DataCache.scala 101:37]
  wire  _GEN_498 = 7'h72 == lineSel ? dirty_114 : _GEN_497; // @[DataCache.scala 101:37]
  wire  _GEN_499 = 7'h73 == lineSel ? dirty_115 : _GEN_498; // @[DataCache.scala 101:37]
  wire  _GEN_500 = 7'h74 == lineSel ? dirty_116 : _GEN_499; // @[DataCache.scala 101:37]
  wire  _GEN_501 = 7'h75 == lineSel ? dirty_117 : _GEN_500; // @[DataCache.scala 101:37]
  wire  _GEN_502 = 7'h76 == lineSel ? dirty_118 : _GEN_501; // @[DataCache.scala 101:37]
  wire  _GEN_503 = 7'h77 == lineSel ? dirty_119 : _GEN_502; // @[DataCache.scala 101:37]
  wire  _GEN_504 = 7'h78 == lineSel ? dirty_120 : _GEN_503; // @[DataCache.scala 101:37]
  wire  _GEN_505 = 7'h79 == lineSel ? dirty_121 : _GEN_504; // @[DataCache.scala 101:37]
  wire  _GEN_506 = 7'h7a == lineSel ? dirty_122 : _GEN_505; // @[DataCache.scala 101:37]
  wire  _GEN_507 = 7'h7b == lineSel ? dirty_123 : _GEN_506; // @[DataCache.scala 101:37]
  wire  _GEN_508 = 7'h7c == lineSel ? dirty_124 : _GEN_507; // @[DataCache.scala 101:37]
  wire  _GEN_509 = 7'h7d == lineSel ? dirty_125 : _GEN_508; // @[DataCache.scala 101:37]
  wire  _GEN_510 = 7'h7e == lineSel ? dirty_126 : _GEN_509; // @[DataCache.scala 101:37]
  wire  _GEN_511 = 7'h7f == lineSel ? dirty_127 : _GEN_510; // @[DataCache.scala 101:37]
  wire  _T_277 = _GEN_127 & _GEN_511; // @[DataCache.scala 101:37]
  wire  _T_278 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_279 = aren & io_axi_readAddr_ready; // @[DataCache.scala 117:18]
  wire  _T_280 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire [4:0] _T_282 = dataOffset + 5'h1; // @[DataCache.scala 126:34]
  wire  _T_283 = io_axi_readData_valid & io_axi_readData_bits_last; // @[DataCache.scala 129:35]
  wire  _GEN_908 = _GEN_3427 | valid_0; // @[DataCache.scala 130:24]
  wire  _GEN_909 = _GEN_3428 | valid_1; // @[DataCache.scala 130:24]
  wire  _GEN_910 = _GEN_3429 | valid_2; // @[DataCache.scala 130:24]
  wire  _GEN_911 = _GEN_3430 | valid_3; // @[DataCache.scala 130:24]
  wire  _GEN_912 = _GEN_3431 | valid_4; // @[DataCache.scala 130:24]
  wire  _GEN_913 = _GEN_3432 | valid_5; // @[DataCache.scala 130:24]
  wire  _GEN_914 = _GEN_3433 | valid_6; // @[DataCache.scala 130:24]
  wire  _GEN_915 = _GEN_3434 | valid_7; // @[DataCache.scala 130:24]
  wire  _GEN_916 = _GEN_3435 | valid_8; // @[DataCache.scala 130:24]
  wire  _GEN_917 = _GEN_3436 | valid_9; // @[DataCache.scala 130:24]
  wire  _GEN_918 = _GEN_3437 | valid_10; // @[DataCache.scala 130:24]
  wire  _GEN_919 = _GEN_3438 | valid_11; // @[DataCache.scala 130:24]
  wire  _GEN_920 = _GEN_3439 | valid_12; // @[DataCache.scala 130:24]
  wire  _GEN_921 = _GEN_3440 | valid_13; // @[DataCache.scala 130:24]
  wire  _GEN_922 = _GEN_3441 | valid_14; // @[DataCache.scala 130:24]
  wire  _GEN_923 = _GEN_3442 | valid_15; // @[DataCache.scala 130:24]
  wire  _GEN_924 = _GEN_3443 | valid_16; // @[DataCache.scala 130:24]
  wire  _GEN_925 = _GEN_3444 | valid_17; // @[DataCache.scala 130:24]
  wire  _GEN_926 = _GEN_3445 | valid_18; // @[DataCache.scala 130:24]
  wire  _GEN_927 = _GEN_3446 | valid_19; // @[DataCache.scala 130:24]
  wire  _GEN_928 = _GEN_3447 | valid_20; // @[DataCache.scala 130:24]
  wire  _GEN_929 = _GEN_3448 | valid_21; // @[DataCache.scala 130:24]
  wire  _GEN_930 = _GEN_3449 | valid_22; // @[DataCache.scala 130:24]
  wire  _GEN_931 = _GEN_3450 | valid_23; // @[DataCache.scala 130:24]
  wire  _GEN_932 = _GEN_3451 | valid_24; // @[DataCache.scala 130:24]
  wire  _GEN_933 = _GEN_3452 | valid_25; // @[DataCache.scala 130:24]
  wire  _GEN_934 = _GEN_3453 | valid_26; // @[DataCache.scala 130:24]
  wire  _GEN_935 = _GEN_3454 | valid_27; // @[DataCache.scala 130:24]
  wire  _GEN_936 = _GEN_3455 | valid_28; // @[DataCache.scala 130:24]
  wire  _GEN_937 = _GEN_3456 | valid_29; // @[DataCache.scala 130:24]
  wire  _GEN_938 = _GEN_3457 | valid_30; // @[DataCache.scala 130:24]
  wire  _GEN_939 = _GEN_3458 | valid_31; // @[DataCache.scala 130:24]
  wire  _GEN_940 = _GEN_3459 | valid_32; // @[DataCache.scala 130:24]
  wire  _GEN_941 = _GEN_3460 | valid_33; // @[DataCache.scala 130:24]
  wire  _GEN_942 = _GEN_3461 | valid_34; // @[DataCache.scala 130:24]
  wire  _GEN_943 = _GEN_3462 | valid_35; // @[DataCache.scala 130:24]
  wire  _GEN_944 = _GEN_3463 | valid_36; // @[DataCache.scala 130:24]
  wire  _GEN_945 = _GEN_3464 | valid_37; // @[DataCache.scala 130:24]
  wire  _GEN_946 = _GEN_3465 | valid_38; // @[DataCache.scala 130:24]
  wire  _GEN_947 = _GEN_3466 | valid_39; // @[DataCache.scala 130:24]
  wire  _GEN_948 = _GEN_3467 | valid_40; // @[DataCache.scala 130:24]
  wire  _GEN_949 = _GEN_3468 | valid_41; // @[DataCache.scala 130:24]
  wire  _GEN_950 = _GEN_3469 | valid_42; // @[DataCache.scala 130:24]
  wire  _GEN_951 = _GEN_3470 | valid_43; // @[DataCache.scala 130:24]
  wire  _GEN_952 = _GEN_3471 | valid_44; // @[DataCache.scala 130:24]
  wire  _GEN_953 = _GEN_3472 | valid_45; // @[DataCache.scala 130:24]
  wire  _GEN_954 = _GEN_3473 | valid_46; // @[DataCache.scala 130:24]
  wire  _GEN_955 = _GEN_3474 | valid_47; // @[DataCache.scala 130:24]
  wire  _GEN_956 = _GEN_3475 | valid_48; // @[DataCache.scala 130:24]
  wire  _GEN_957 = _GEN_3476 | valid_49; // @[DataCache.scala 130:24]
  wire  _GEN_958 = _GEN_3477 | valid_50; // @[DataCache.scala 130:24]
  wire  _GEN_959 = _GEN_3478 | valid_51; // @[DataCache.scala 130:24]
  wire  _GEN_960 = _GEN_3479 | valid_52; // @[DataCache.scala 130:24]
  wire  _GEN_961 = _GEN_3480 | valid_53; // @[DataCache.scala 130:24]
  wire  _GEN_962 = _GEN_3481 | valid_54; // @[DataCache.scala 130:24]
  wire  _GEN_963 = _GEN_3482 | valid_55; // @[DataCache.scala 130:24]
  wire  _GEN_964 = _GEN_3483 | valid_56; // @[DataCache.scala 130:24]
  wire  _GEN_965 = _GEN_3484 | valid_57; // @[DataCache.scala 130:24]
  wire  _GEN_966 = _GEN_3485 | valid_58; // @[DataCache.scala 130:24]
  wire  _GEN_967 = _GEN_3486 | valid_59; // @[DataCache.scala 130:24]
  wire  _GEN_968 = _GEN_3487 | valid_60; // @[DataCache.scala 130:24]
  wire  _GEN_969 = _GEN_3488 | valid_61; // @[DataCache.scala 130:24]
  wire  _GEN_970 = _GEN_3489 | valid_62; // @[DataCache.scala 130:24]
  wire  _GEN_971 = _GEN_3490 | valid_63; // @[DataCache.scala 130:24]
  wire  _GEN_972 = _GEN_3491 | valid_64; // @[DataCache.scala 130:24]
  wire  _GEN_973 = _GEN_3492 | valid_65; // @[DataCache.scala 130:24]
  wire  _GEN_974 = _GEN_3493 | valid_66; // @[DataCache.scala 130:24]
  wire  _GEN_975 = _GEN_3494 | valid_67; // @[DataCache.scala 130:24]
  wire  _GEN_976 = _GEN_3495 | valid_68; // @[DataCache.scala 130:24]
  wire  _GEN_977 = _GEN_3496 | valid_69; // @[DataCache.scala 130:24]
  wire  _GEN_978 = _GEN_3497 | valid_70; // @[DataCache.scala 130:24]
  wire  _GEN_979 = _GEN_3498 | valid_71; // @[DataCache.scala 130:24]
  wire  _GEN_980 = _GEN_3499 | valid_72; // @[DataCache.scala 130:24]
  wire  _GEN_981 = _GEN_3500 | valid_73; // @[DataCache.scala 130:24]
  wire  _GEN_982 = _GEN_3501 | valid_74; // @[DataCache.scala 130:24]
  wire  _GEN_983 = _GEN_3502 | valid_75; // @[DataCache.scala 130:24]
  wire  _GEN_984 = _GEN_3503 | valid_76; // @[DataCache.scala 130:24]
  wire  _GEN_985 = _GEN_3504 | valid_77; // @[DataCache.scala 130:24]
  wire  _GEN_986 = _GEN_3505 | valid_78; // @[DataCache.scala 130:24]
  wire  _GEN_987 = _GEN_3506 | valid_79; // @[DataCache.scala 130:24]
  wire  _GEN_988 = _GEN_3507 | valid_80; // @[DataCache.scala 130:24]
  wire  _GEN_989 = _GEN_3508 | valid_81; // @[DataCache.scala 130:24]
  wire  _GEN_990 = _GEN_3509 | valid_82; // @[DataCache.scala 130:24]
  wire  _GEN_991 = _GEN_3510 | valid_83; // @[DataCache.scala 130:24]
  wire  _GEN_992 = _GEN_3511 | valid_84; // @[DataCache.scala 130:24]
  wire  _GEN_993 = _GEN_3512 | valid_85; // @[DataCache.scala 130:24]
  wire  _GEN_994 = _GEN_3513 | valid_86; // @[DataCache.scala 130:24]
  wire  _GEN_995 = _GEN_3514 | valid_87; // @[DataCache.scala 130:24]
  wire  _GEN_996 = _GEN_3515 | valid_88; // @[DataCache.scala 130:24]
  wire  _GEN_997 = _GEN_3516 | valid_89; // @[DataCache.scala 130:24]
  wire  _GEN_998 = _GEN_3517 | valid_90; // @[DataCache.scala 130:24]
  wire  _GEN_999 = _GEN_3518 | valid_91; // @[DataCache.scala 130:24]
  wire  _GEN_1000 = _GEN_3519 | valid_92; // @[DataCache.scala 130:24]
  wire  _GEN_1001 = _GEN_3520 | valid_93; // @[DataCache.scala 130:24]
  wire  _GEN_1002 = _GEN_3521 | valid_94; // @[DataCache.scala 130:24]
  wire  _GEN_1003 = _GEN_3522 | valid_95; // @[DataCache.scala 130:24]
  wire  _GEN_1004 = _GEN_3523 | valid_96; // @[DataCache.scala 130:24]
  wire  _GEN_1005 = _GEN_3524 | valid_97; // @[DataCache.scala 130:24]
  wire  _GEN_1006 = _GEN_3525 | valid_98; // @[DataCache.scala 130:24]
  wire  _GEN_1007 = _GEN_3526 | valid_99; // @[DataCache.scala 130:24]
  wire  _GEN_1008 = _GEN_3527 | valid_100; // @[DataCache.scala 130:24]
  wire  _GEN_1009 = _GEN_3528 | valid_101; // @[DataCache.scala 130:24]
  wire  _GEN_1010 = _GEN_3529 | valid_102; // @[DataCache.scala 130:24]
  wire  _GEN_1011 = _GEN_3530 | valid_103; // @[DataCache.scala 130:24]
  wire  _GEN_1012 = _GEN_3531 | valid_104; // @[DataCache.scala 130:24]
  wire  _GEN_1013 = _GEN_3532 | valid_105; // @[DataCache.scala 130:24]
  wire  _GEN_1014 = _GEN_3533 | valid_106; // @[DataCache.scala 130:24]
  wire  _GEN_1015 = _GEN_3534 | valid_107; // @[DataCache.scala 130:24]
  wire  _GEN_1016 = _GEN_3535 | valid_108; // @[DataCache.scala 130:24]
  wire  _GEN_1017 = _GEN_3536 | valid_109; // @[DataCache.scala 130:24]
  wire  _GEN_1018 = _GEN_3537 | valid_110; // @[DataCache.scala 130:24]
  wire  _GEN_1019 = _GEN_3538 | valid_111; // @[DataCache.scala 130:24]
  wire  _GEN_1020 = _GEN_3539 | valid_112; // @[DataCache.scala 130:24]
  wire  _GEN_1021 = _GEN_3540 | valid_113; // @[DataCache.scala 130:24]
  wire  _GEN_1022 = _GEN_3541 | valid_114; // @[DataCache.scala 130:24]
  wire  _GEN_1023 = _GEN_3542 | valid_115; // @[DataCache.scala 130:24]
  wire  _GEN_1024 = _GEN_3543 | valid_116; // @[DataCache.scala 130:24]
  wire  _GEN_1025 = _GEN_3544 | valid_117; // @[DataCache.scala 130:24]
  wire  _GEN_1026 = _GEN_3545 | valid_118; // @[DataCache.scala 130:24]
  wire  _GEN_1027 = _GEN_3546 | valid_119; // @[DataCache.scala 130:24]
  wire  _GEN_1028 = _GEN_3547 | valid_120; // @[DataCache.scala 130:24]
  wire  _GEN_1029 = _GEN_3548 | valid_121; // @[DataCache.scala 130:24]
  wire  _GEN_1030 = _GEN_3549 | valid_122; // @[DataCache.scala 130:24]
  wire  _GEN_1031 = _GEN_3550 | valid_123; // @[DataCache.scala 130:24]
  wire  _GEN_1032 = _GEN_3551 | valid_124; // @[DataCache.scala 130:24]
  wire  _GEN_1033 = _GEN_3552 | valid_125; // @[DataCache.scala 130:24]
  wire  _GEN_1034 = _GEN_3553 | valid_126; // @[DataCache.scala 130:24]
  wire  _GEN_1035 = _GEN_3554 | valid_127; // @[DataCache.scala 130:24]
  wire  _T_285 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_286 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_287 = awen & io_axi_writeAddr_ready; // @[DataCache.scala 145:18]
  wire  _T_288 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_289 = ~wlast; // @[DataCache.scala 155:39]
  wire  _T_290 = io_axi_writeData_ready & _T_289; // @[DataCache.scala 155:36]
  wire  _T_293 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_295 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire  _T_300 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire  _GEN_2880 = _T_280 & _T_283; // @[Conditional.scala 39:67]
  wire  _GEN_3150 = _T_278 ? 1'h0 : _GEN_2880; // @[Conditional.scala 39:67]
  wire  _T_303 = ~isDirty; // @[DataCache.scala 204:53]
  wire  _T_304 = io_flush ? _T_303 : cacheHit; // @[DataCache.scala 204:42]
  BlockMem lines ( // @[DataCache.scala 40:21]
    .clock(lines_clock),
    .io_wen(lines_io_wen),
    .io_addr(lines_io_addr),
    .io_wdata(lines_io_wdata),
    .io_rdata(lines_io_rdata)
  );
  assign tag__T_4_addr = selAddr[12:6];
  assign tag__T_4_data = tag[tag__T_4_addr]; // @[DataCache.scala 39:18]
  assign tag__T_6_addr = selAddr[12:6];
  assign tag__T_6_data = tag[tag__T_6_addr]; // @[DataCache.scala 39:18]
  assign tag__T_261_addr = realDirty_0 ? 7'h0 : _T_259;
  assign tag__T_261_data = tag[tag__T_261_addr]; // @[DataCache.scala 39:18]
  assign tag__T_284_data = selAddr[31:13];
  assign tag__T_284_addr = selAddr[12:6];
  assign tag__T_284_mask = 1'h1;
  assign tag__T_284_en = _T_274 ? 1'h0 : _GEN_3150;
  assign io_sram_valid = _T_2 & _T_304; // @[DataCache.scala 204:17]
  assign io_sram_rdata = lines_io_rdata; // @[DataCache.scala 206:17]
  assign io_axi_readAddr_valid = aren; // @[AXI.scala 56:20 DataCache.scala 210:31]
  assign io_axi_readAddr_bits_addr = raddr; // @[AXI.scala 9:21 DataCache.scala 211:31]
  assign io_axi_writeAddr_valid = awen; // @[AXI.scala 59:21 DataCache.scala 216:31]
  assign io_axi_writeAddr_bits_addr = waddr; // @[AXI.scala 9:21 DataCache.scala 217:31]
  assign io_axi_writeData_valid = wen; // @[AXI.scala 61:21 DataCache.scala 221:31]
  assign io_axi_writeData_bits_data = lines_io_rdata; // @[AXI.scala 9:21 DataCache.scala 222:31]
  assign io_axi_writeData_bits_last = wen & _T_1; // @[AXI.scala 9:21 DataCache.scala 223:31]
  assign lines_clock = clock;
  assign lines_io_wen = lineEnCpu ? io_sram_wen : _T_268; // @[DataCache.scala 80:19]
  assign lines_io_addr = _T_270 ? dataSel : _T_271; // @[DataCache.scala 82:19]
  assign lines_io_wdata = lineEnCpu ? io_sram_wdata : io_axi_readData_bits_data; // @[DataCache.scala 84:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    tag[initvar] = _RAND_0[18:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  valid_0 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  valid_1 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  valid_2 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  valid_3 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  valid_4 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  valid_5 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  valid_6 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  valid_7 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  valid_8 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  valid_9 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  valid_10 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  valid_11 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  valid_12 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  valid_13 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  valid_14 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  valid_15 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  valid_16 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  valid_17 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  valid_18 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  valid_19 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  valid_20 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  valid_21 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  valid_22 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  valid_23 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  valid_24 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  valid_25 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  valid_26 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  valid_27 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  valid_28 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  valid_29 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  valid_30 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  valid_31 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  valid_32 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  valid_33 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  valid_34 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  valid_35 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  valid_36 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  valid_37 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  valid_38 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  valid_39 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  valid_40 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  valid_41 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  valid_42 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  valid_43 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  valid_44 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  valid_45 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  valid_46 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  valid_47 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  valid_48 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  valid_49 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  valid_50 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  valid_51 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  valid_52 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  valid_53 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  valid_54 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  valid_55 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  valid_56 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  valid_57 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  valid_58 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  valid_59 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  valid_60 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  valid_61 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  valid_62 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  valid_63 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  valid_64 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  valid_65 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  valid_66 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  valid_67 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  valid_68 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  valid_69 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  valid_70 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  valid_71 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  valid_72 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  valid_73 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  valid_74 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  valid_75 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  valid_76 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  valid_77 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  valid_78 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  valid_79 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  valid_80 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  valid_81 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  valid_82 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  valid_83 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  valid_84 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  valid_85 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  valid_86 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  valid_87 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  valid_88 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  valid_89 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  valid_90 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  valid_91 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  valid_92 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  valid_93 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  valid_94 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  valid_95 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  valid_96 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  valid_97 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  valid_98 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  valid_99 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  valid_100 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  valid_101 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  valid_102 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  valid_103 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  valid_104 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  valid_105 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  valid_106 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  valid_107 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  valid_108 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  valid_109 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  valid_110 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  valid_111 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  valid_112 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  valid_113 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  valid_114 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  valid_115 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  valid_116 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  valid_117 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  valid_118 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  valid_119 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  valid_120 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  valid_121 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  valid_122 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  valid_123 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  valid_124 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  valid_125 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  valid_126 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  valid_127 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  dirty_0 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  dirty_1 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  dirty_2 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  dirty_3 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  dirty_4 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  dirty_5 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  dirty_6 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  dirty_7 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  dirty_8 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  dirty_9 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  dirty_10 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  dirty_11 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  dirty_12 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  dirty_13 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  dirty_14 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  dirty_15 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  dirty_16 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  dirty_17 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  dirty_18 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  dirty_19 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  dirty_20 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  dirty_21 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  dirty_22 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  dirty_23 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  dirty_24 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  dirty_25 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  dirty_26 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  dirty_27 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  dirty_28 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  dirty_29 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  dirty_30 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  dirty_31 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  dirty_32 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  dirty_33 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  dirty_34 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  dirty_35 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  dirty_36 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  dirty_37 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  dirty_38 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  dirty_39 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  dirty_40 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  dirty_41 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  dirty_42 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  dirty_43 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  dirty_44 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  dirty_45 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  dirty_46 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  dirty_47 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  dirty_48 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  dirty_49 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  dirty_50 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  dirty_51 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  dirty_52 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  dirty_53 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  dirty_54 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  dirty_55 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  dirty_56 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  dirty_57 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  dirty_58 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  dirty_59 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  dirty_60 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  dirty_61 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  dirty_62 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  dirty_63 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  dirty_64 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  dirty_65 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  dirty_66 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  dirty_67 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  dirty_68 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  dirty_69 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  dirty_70 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  dirty_71 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  dirty_72 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  dirty_73 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  dirty_74 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  dirty_75 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  dirty_76 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  dirty_77 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  dirty_78 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  dirty_79 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  dirty_80 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  dirty_81 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  dirty_82 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  dirty_83 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  dirty_84 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  dirty_85 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  dirty_86 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  dirty_87 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  dirty_88 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  dirty_89 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  dirty_90 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  dirty_91 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  dirty_92 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  dirty_93 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  dirty_94 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  dirty_95 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  dirty_96 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  dirty_97 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  dirty_98 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  dirty_99 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  dirty_100 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  dirty_101 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  dirty_102 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  dirty_103 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  dirty_104 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  dirty_105 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  dirty_106 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  dirty_107 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  dirty_108 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  dirty_109 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  dirty_110 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  dirty_111 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  dirty_112 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  dirty_113 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  dirty_114 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  dirty_115 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  dirty_116 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  dirty_117 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  dirty_118 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  dirty_119 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  dirty_120 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  dirty_121 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  dirty_122 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  dirty_123 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  dirty_124 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  dirty_125 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  dirty_126 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  dirty_127 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  dataOffset = _RAND_258[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  lastOffset = _RAND_259[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  aren = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  raddr = _RAND_261[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  awen = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  waddr = _RAND_263[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  wen = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  sramAddr = _RAND_265[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tag__T_284_en & tag__T_284_mask) begin
      tag[tag__T_284_addr] <= tag__T_284_data; // @[DataCache.scala 39:18]
    end
    if (reset) begin
      state <= 4'h0;
    end else if (_T_274) begin
      if (_T_275) begin
        state <= 4'h6;
      end else if (io_sram_en) begin
        if (!(cacheHit)) begin
          if (_T_277) begin
            state <= 4'h4;
          end else begin
            state <= 4'h1;
          end
        end
      end
    end else if (_T_278) begin
      if (_T_279) begin
        state <= 4'h2;
      end
    end else if (_T_280) begin
      if (_T_283) begin
        state <= 4'h3;
      end
    end else if (_T_285) begin
      state <= 4'h0;
    end else if (_T_286) begin
      if (_T_287) begin
        state <= 4'h5;
      end
    end else if (_T_288) begin
      if (wlast) begin
        state <= 4'h1;
      end
    end else if (_T_293) begin
      if (_T_287) begin
        state <= 4'h7;
      end
    end else if (_T_295) begin
      if (wlast) begin
        state <= 4'h8;
      end
    end else if (_T_300) begin
      if (isDirty) begin
        state <= 4'h6;
      end else begin
        state <= 4'h0;
      end
    end
    if (reset) begin
      valid_0 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_0 <= _GEN_908;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h0 == lineSel) begin
                  valid_0 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h0 == nextDirty) begin
                    valid_0 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_1 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_1 <= _GEN_909;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h1 == lineSel) begin
                  valid_1 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h1 == nextDirty) begin
                    valid_1 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_2 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_2 <= _GEN_910;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h2 == lineSel) begin
                  valid_2 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h2 == nextDirty) begin
                    valid_2 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_3 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_3 <= _GEN_911;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h3 == lineSel) begin
                  valid_3 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h3 == nextDirty) begin
                    valid_3 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_4 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_4 <= _GEN_912;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h4 == lineSel) begin
                  valid_4 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h4 == nextDirty) begin
                    valid_4 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_5 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_5 <= _GEN_913;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h5 == lineSel) begin
                  valid_5 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h5 == nextDirty) begin
                    valid_5 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_6 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_6 <= _GEN_914;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h6 == lineSel) begin
                  valid_6 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h6 == nextDirty) begin
                    valid_6 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_7 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_7 <= _GEN_915;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h7 == lineSel) begin
                  valid_7 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h7 == nextDirty) begin
                    valid_7 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_8 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_8 <= _GEN_916;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h8 == lineSel) begin
                  valid_8 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h8 == nextDirty) begin
                    valid_8 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_9 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_9 <= _GEN_917;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h9 == lineSel) begin
                  valid_9 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h9 == nextDirty) begin
                    valid_9 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_10 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_10 <= _GEN_918;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'ha == lineSel) begin
                  valid_10 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'ha == nextDirty) begin
                    valid_10 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_11 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_11 <= _GEN_919;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'hb == lineSel) begin
                  valid_11 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'hb == nextDirty) begin
                    valid_11 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_12 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_12 <= _GEN_920;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'hc == lineSel) begin
                  valid_12 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'hc == nextDirty) begin
                    valid_12 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_13 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_13 <= _GEN_921;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'hd == lineSel) begin
                  valid_13 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'hd == nextDirty) begin
                    valid_13 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_14 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_14 <= _GEN_922;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'he == lineSel) begin
                  valid_14 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'he == nextDirty) begin
                    valid_14 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_15 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_15 <= _GEN_923;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'hf == lineSel) begin
                  valid_15 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'hf == nextDirty) begin
                    valid_15 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_16 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_16 <= _GEN_924;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h10 == lineSel) begin
                  valid_16 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h10 == nextDirty) begin
                    valid_16 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_17 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_17 <= _GEN_925;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h11 == lineSel) begin
                  valid_17 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h11 == nextDirty) begin
                    valid_17 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_18 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_18 <= _GEN_926;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h12 == lineSel) begin
                  valid_18 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h12 == nextDirty) begin
                    valid_18 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_19 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_19 <= _GEN_927;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h13 == lineSel) begin
                  valid_19 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h13 == nextDirty) begin
                    valid_19 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_20 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_20 <= _GEN_928;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h14 == lineSel) begin
                  valid_20 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h14 == nextDirty) begin
                    valid_20 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_21 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_21 <= _GEN_929;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h15 == lineSel) begin
                  valid_21 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h15 == nextDirty) begin
                    valid_21 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_22 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_22 <= _GEN_930;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h16 == lineSel) begin
                  valid_22 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h16 == nextDirty) begin
                    valid_22 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_23 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_23 <= _GEN_931;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h17 == lineSel) begin
                  valid_23 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h17 == nextDirty) begin
                    valid_23 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_24 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_24 <= _GEN_932;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h18 == lineSel) begin
                  valid_24 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h18 == nextDirty) begin
                    valid_24 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_25 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_25 <= _GEN_933;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h19 == lineSel) begin
                  valid_25 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h19 == nextDirty) begin
                    valid_25 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_26 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_26 <= _GEN_934;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h1a == lineSel) begin
                  valid_26 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h1a == nextDirty) begin
                    valid_26 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_27 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_27 <= _GEN_935;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h1b == lineSel) begin
                  valid_27 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h1b == nextDirty) begin
                    valid_27 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_28 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_28 <= _GEN_936;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h1c == lineSel) begin
                  valid_28 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h1c == nextDirty) begin
                    valid_28 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_29 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_29 <= _GEN_937;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h1d == lineSel) begin
                  valid_29 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h1d == nextDirty) begin
                    valid_29 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_30 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_30 <= _GEN_938;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h1e == lineSel) begin
                  valid_30 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h1e == nextDirty) begin
                    valid_30 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_31 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_31 <= _GEN_939;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h1f == lineSel) begin
                  valid_31 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h1f == nextDirty) begin
                    valid_31 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_32 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_32 <= _GEN_940;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h20 == lineSel) begin
                  valid_32 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h20 == nextDirty) begin
                    valid_32 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_33 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_33 <= _GEN_941;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h21 == lineSel) begin
                  valid_33 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h21 == nextDirty) begin
                    valid_33 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_34 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_34 <= _GEN_942;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h22 == lineSel) begin
                  valid_34 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h22 == nextDirty) begin
                    valid_34 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_35 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_35 <= _GEN_943;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h23 == lineSel) begin
                  valid_35 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h23 == nextDirty) begin
                    valid_35 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_36 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_36 <= _GEN_944;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h24 == lineSel) begin
                  valid_36 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h24 == nextDirty) begin
                    valid_36 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_37 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_37 <= _GEN_945;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h25 == lineSel) begin
                  valid_37 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h25 == nextDirty) begin
                    valid_37 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_38 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_38 <= _GEN_946;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h26 == lineSel) begin
                  valid_38 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h26 == nextDirty) begin
                    valid_38 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_39 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_39 <= _GEN_947;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h27 == lineSel) begin
                  valid_39 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h27 == nextDirty) begin
                    valid_39 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_40 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_40 <= _GEN_948;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h28 == lineSel) begin
                  valid_40 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h28 == nextDirty) begin
                    valid_40 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_41 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_41 <= _GEN_949;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h29 == lineSel) begin
                  valid_41 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h29 == nextDirty) begin
                    valid_41 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_42 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_42 <= _GEN_950;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h2a == lineSel) begin
                  valid_42 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h2a == nextDirty) begin
                    valid_42 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_43 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_43 <= _GEN_951;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h2b == lineSel) begin
                  valid_43 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h2b == nextDirty) begin
                    valid_43 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_44 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_44 <= _GEN_952;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h2c == lineSel) begin
                  valid_44 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h2c == nextDirty) begin
                    valid_44 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_45 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_45 <= _GEN_953;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h2d == lineSel) begin
                  valid_45 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h2d == nextDirty) begin
                    valid_45 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_46 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_46 <= _GEN_954;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h2e == lineSel) begin
                  valid_46 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h2e == nextDirty) begin
                    valid_46 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_47 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_47 <= _GEN_955;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h2f == lineSel) begin
                  valid_47 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h2f == nextDirty) begin
                    valid_47 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_48 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_48 <= _GEN_956;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h30 == lineSel) begin
                  valid_48 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h30 == nextDirty) begin
                    valid_48 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_49 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_49 <= _GEN_957;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h31 == lineSel) begin
                  valid_49 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h31 == nextDirty) begin
                    valid_49 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_50 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_50 <= _GEN_958;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h32 == lineSel) begin
                  valid_50 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h32 == nextDirty) begin
                    valid_50 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_51 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_51 <= _GEN_959;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h33 == lineSel) begin
                  valid_51 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h33 == nextDirty) begin
                    valid_51 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_52 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_52 <= _GEN_960;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h34 == lineSel) begin
                  valid_52 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h34 == nextDirty) begin
                    valid_52 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_53 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_53 <= _GEN_961;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h35 == lineSel) begin
                  valid_53 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h35 == nextDirty) begin
                    valid_53 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_54 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_54 <= _GEN_962;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h36 == lineSel) begin
                  valid_54 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h36 == nextDirty) begin
                    valid_54 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_55 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_55 <= _GEN_963;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h37 == lineSel) begin
                  valid_55 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h37 == nextDirty) begin
                    valid_55 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_56 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_56 <= _GEN_964;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h38 == lineSel) begin
                  valid_56 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h38 == nextDirty) begin
                    valid_56 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_57 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_57 <= _GEN_965;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h39 == lineSel) begin
                  valid_57 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h39 == nextDirty) begin
                    valid_57 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_58 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_58 <= _GEN_966;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h3a == lineSel) begin
                  valid_58 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h3a == nextDirty) begin
                    valid_58 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_59 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_59 <= _GEN_967;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h3b == lineSel) begin
                  valid_59 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h3b == nextDirty) begin
                    valid_59 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_60 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_60 <= _GEN_968;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h3c == lineSel) begin
                  valid_60 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h3c == nextDirty) begin
                    valid_60 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_61 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_61 <= _GEN_969;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h3d == lineSel) begin
                  valid_61 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h3d == nextDirty) begin
                    valid_61 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_62 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_62 <= _GEN_970;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h3e == lineSel) begin
                  valid_62 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h3e == nextDirty) begin
                    valid_62 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_63 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_63 <= _GEN_971;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h3f == lineSel) begin
                  valid_63 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h3f == nextDirty) begin
                    valid_63 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_64 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_64 <= _GEN_972;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h40 == lineSel) begin
                  valid_64 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h40 == nextDirty) begin
                    valid_64 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_65 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_65 <= _GEN_973;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h41 == lineSel) begin
                  valid_65 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h41 == nextDirty) begin
                    valid_65 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_66 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_66 <= _GEN_974;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h42 == lineSel) begin
                  valid_66 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h42 == nextDirty) begin
                    valid_66 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_67 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_67 <= _GEN_975;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h43 == lineSel) begin
                  valid_67 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h43 == nextDirty) begin
                    valid_67 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_68 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_68 <= _GEN_976;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h44 == lineSel) begin
                  valid_68 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h44 == nextDirty) begin
                    valid_68 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_69 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_69 <= _GEN_977;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h45 == lineSel) begin
                  valid_69 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h45 == nextDirty) begin
                    valid_69 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_70 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_70 <= _GEN_978;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h46 == lineSel) begin
                  valid_70 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h46 == nextDirty) begin
                    valid_70 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_71 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_71 <= _GEN_979;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h47 == lineSel) begin
                  valid_71 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h47 == nextDirty) begin
                    valid_71 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_72 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_72 <= _GEN_980;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h48 == lineSel) begin
                  valid_72 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h48 == nextDirty) begin
                    valid_72 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_73 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_73 <= _GEN_981;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h49 == lineSel) begin
                  valid_73 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h49 == nextDirty) begin
                    valid_73 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_74 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_74 <= _GEN_982;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h4a == lineSel) begin
                  valid_74 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h4a == nextDirty) begin
                    valid_74 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_75 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_75 <= _GEN_983;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h4b == lineSel) begin
                  valid_75 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h4b == nextDirty) begin
                    valid_75 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_76 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_76 <= _GEN_984;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h4c == lineSel) begin
                  valid_76 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h4c == nextDirty) begin
                    valid_76 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_77 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_77 <= _GEN_985;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h4d == lineSel) begin
                  valid_77 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h4d == nextDirty) begin
                    valid_77 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_78 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_78 <= _GEN_986;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h4e == lineSel) begin
                  valid_78 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h4e == nextDirty) begin
                    valid_78 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_79 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_79 <= _GEN_987;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h4f == lineSel) begin
                  valid_79 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h4f == nextDirty) begin
                    valid_79 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_80 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_80 <= _GEN_988;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h50 == lineSel) begin
                  valid_80 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h50 == nextDirty) begin
                    valid_80 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_81 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_81 <= _GEN_989;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h51 == lineSel) begin
                  valid_81 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h51 == nextDirty) begin
                    valid_81 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_82 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_82 <= _GEN_990;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h52 == lineSel) begin
                  valid_82 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h52 == nextDirty) begin
                    valid_82 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_83 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_83 <= _GEN_991;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h53 == lineSel) begin
                  valid_83 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h53 == nextDirty) begin
                    valid_83 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_84 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_84 <= _GEN_992;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h54 == lineSel) begin
                  valid_84 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h54 == nextDirty) begin
                    valid_84 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_85 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_85 <= _GEN_993;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h55 == lineSel) begin
                  valid_85 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h55 == nextDirty) begin
                    valid_85 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_86 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_86 <= _GEN_994;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h56 == lineSel) begin
                  valid_86 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h56 == nextDirty) begin
                    valid_86 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_87 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_87 <= _GEN_995;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h57 == lineSel) begin
                  valid_87 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h57 == nextDirty) begin
                    valid_87 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_88 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_88 <= _GEN_996;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h58 == lineSel) begin
                  valid_88 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h58 == nextDirty) begin
                    valid_88 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_89 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_89 <= _GEN_997;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h59 == lineSel) begin
                  valid_89 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h59 == nextDirty) begin
                    valid_89 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_90 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_90 <= _GEN_998;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h5a == lineSel) begin
                  valid_90 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h5a == nextDirty) begin
                    valid_90 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_91 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_91 <= _GEN_999;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h5b == lineSel) begin
                  valid_91 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h5b == nextDirty) begin
                    valid_91 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_92 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_92 <= _GEN_1000;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h5c == lineSel) begin
                  valid_92 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h5c == nextDirty) begin
                    valid_92 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_93 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_93 <= _GEN_1001;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h5d == lineSel) begin
                  valid_93 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h5d == nextDirty) begin
                    valid_93 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_94 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_94 <= _GEN_1002;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h5e == lineSel) begin
                  valid_94 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h5e == nextDirty) begin
                    valid_94 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_95 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_95 <= _GEN_1003;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h5f == lineSel) begin
                  valid_95 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h5f == nextDirty) begin
                    valid_95 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_96 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_96 <= _GEN_1004;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h60 == lineSel) begin
                  valid_96 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h60 == nextDirty) begin
                    valid_96 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_97 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_97 <= _GEN_1005;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h61 == lineSel) begin
                  valid_97 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h61 == nextDirty) begin
                    valid_97 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_98 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_98 <= _GEN_1006;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h62 == lineSel) begin
                  valid_98 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h62 == nextDirty) begin
                    valid_98 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_99 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_99 <= _GEN_1007;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h63 == lineSel) begin
                  valid_99 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h63 == nextDirty) begin
                    valid_99 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_100 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_100 <= _GEN_1008;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h64 == lineSel) begin
                  valid_100 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h64 == nextDirty) begin
                    valid_100 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_101 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_101 <= _GEN_1009;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h65 == lineSel) begin
                  valid_101 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h65 == nextDirty) begin
                    valid_101 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_102 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_102 <= _GEN_1010;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h66 == lineSel) begin
                  valid_102 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h66 == nextDirty) begin
                    valid_102 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_103 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_103 <= _GEN_1011;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h67 == lineSel) begin
                  valid_103 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h67 == nextDirty) begin
                    valid_103 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_104 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_104 <= _GEN_1012;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h68 == lineSel) begin
                  valid_104 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h68 == nextDirty) begin
                    valid_104 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_105 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_105 <= _GEN_1013;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h69 == lineSel) begin
                  valid_105 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h69 == nextDirty) begin
                    valid_105 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_106 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_106 <= _GEN_1014;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h6a == lineSel) begin
                  valid_106 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h6a == nextDirty) begin
                    valid_106 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_107 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_107 <= _GEN_1015;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h6b == lineSel) begin
                  valid_107 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h6b == nextDirty) begin
                    valid_107 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_108 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_108 <= _GEN_1016;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h6c == lineSel) begin
                  valid_108 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h6c == nextDirty) begin
                    valid_108 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_109 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_109 <= _GEN_1017;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h6d == lineSel) begin
                  valid_109 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h6d == nextDirty) begin
                    valid_109 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_110 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_110 <= _GEN_1018;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h6e == lineSel) begin
                  valid_110 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h6e == nextDirty) begin
                    valid_110 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_111 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_111 <= _GEN_1019;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h6f == lineSel) begin
                  valid_111 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h6f == nextDirty) begin
                    valid_111 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_112 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_112 <= _GEN_1020;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h70 == lineSel) begin
                  valid_112 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h70 == nextDirty) begin
                    valid_112 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_113 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_113 <= _GEN_1021;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h71 == lineSel) begin
                  valid_113 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h71 == nextDirty) begin
                    valid_113 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_114 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_114 <= _GEN_1022;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h72 == lineSel) begin
                  valid_114 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h72 == nextDirty) begin
                    valid_114 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_115 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_115 <= _GEN_1023;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h73 == lineSel) begin
                  valid_115 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h73 == nextDirty) begin
                    valid_115 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_116 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_116 <= _GEN_1024;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h74 == lineSel) begin
                  valid_116 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h74 == nextDirty) begin
                    valid_116 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_117 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_117 <= _GEN_1025;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h75 == lineSel) begin
                  valid_117 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h75 == nextDirty) begin
                    valid_117 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_118 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_118 <= _GEN_1026;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h76 == lineSel) begin
                  valid_118 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h76 == nextDirty) begin
                    valid_118 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_119 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_119 <= _GEN_1027;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h77 == lineSel) begin
                  valid_119 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h77 == nextDirty) begin
                    valid_119 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_120 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_120 <= _GEN_1028;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h78 == lineSel) begin
                  valid_120 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h78 == nextDirty) begin
                    valid_120 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_121 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_121 <= _GEN_1029;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h79 == lineSel) begin
                  valid_121 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h79 == nextDirty) begin
                    valid_121 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_122 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_122 <= _GEN_1030;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h7a == lineSel) begin
                  valid_122 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h7a == nextDirty) begin
                    valid_122 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_123 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_123 <= _GEN_1031;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h7b == lineSel) begin
                  valid_123 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h7b == nextDirty) begin
                    valid_123 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_124 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_124 <= _GEN_1032;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h7c == lineSel) begin
                  valid_124 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h7c == nextDirty) begin
                    valid_124 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_125 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_125 <= _GEN_1033;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h7d == lineSel) begin
                  valid_125 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h7d == nextDirty) begin
                    valid_125 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_126 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_126 <= _GEN_1034;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h7e == lineSel) begin
                  valid_126 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h7e == nextDirty) begin
                    valid_126 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      valid_127 <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (_T_280) begin
          if (_T_283) begin
            valid_127 <= _GEN_1035;
          end
        end else if (!(_T_285)) begin
          if (!(_T_286)) begin
            if (_T_288) begin
              if (wlast) begin
                if (7'h7f == lineSel) begin
                  valid_127 <= 1'h0;
                end
              end
            end else if (!(_T_293)) begin
              if (_T_295) begin
                if (wlast) begin
                  if (7'h7f == nextDirty) begin
                    valid_127 <= 1'h0;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_0 <= _GEN_128;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h0 == lineSel) begin
            dirty_0 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_1 <= _GEN_129;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h1 == lineSel) begin
            dirty_1 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_2 <= _GEN_130;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h2 == lineSel) begin
            dirty_2 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_3 <= _GEN_131;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h3 == lineSel) begin
            dirty_3 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_4 <= _GEN_132;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h4 == lineSel) begin
            dirty_4 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_5 <= _GEN_133;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h5 == lineSel) begin
            dirty_5 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_6 <= _GEN_134;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h6 == lineSel) begin
            dirty_6 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_7 <= _GEN_135;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h7 == lineSel) begin
            dirty_7 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_8 <= _GEN_136;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h8 == lineSel) begin
            dirty_8 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_9 <= _GEN_137;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h9 == lineSel) begin
            dirty_9 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_10 <= _GEN_138;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'ha == lineSel) begin
            dirty_10 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_11 <= _GEN_139;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'hb == lineSel) begin
            dirty_11 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_12 <= _GEN_140;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'hc == lineSel) begin
            dirty_12 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_13 <= _GEN_141;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'hd == lineSel) begin
            dirty_13 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_14 <= _GEN_142;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'he == lineSel) begin
            dirty_14 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_15 <= _GEN_143;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'hf == lineSel) begin
            dirty_15 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_16 <= _GEN_144;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h10 == lineSel) begin
            dirty_16 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_17 <= _GEN_145;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h11 == lineSel) begin
            dirty_17 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_18 <= _GEN_146;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h12 == lineSel) begin
            dirty_18 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_19 <= _GEN_147;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h13 == lineSel) begin
            dirty_19 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_20 <= _GEN_148;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h14 == lineSel) begin
            dirty_20 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_21 <= _GEN_149;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h15 == lineSel) begin
            dirty_21 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_22 <= _GEN_150;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h16 == lineSel) begin
            dirty_22 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_23 <= _GEN_151;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h17 == lineSel) begin
            dirty_23 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_24 <= _GEN_152;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h18 == lineSel) begin
            dirty_24 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_25 <= _GEN_153;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h19 == lineSel) begin
            dirty_25 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_26 <= _GEN_154;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h1a == lineSel) begin
            dirty_26 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_27 <= _GEN_155;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h1b == lineSel) begin
            dirty_27 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_28 <= _GEN_156;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h1c == lineSel) begin
            dirty_28 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_29 <= _GEN_157;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h1d == lineSel) begin
            dirty_29 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_30 <= _GEN_158;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h1e == lineSel) begin
            dirty_30 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_31 <= _GEN_159;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h1f == lineSel) begin
            dirty_31 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_32 <= _GEN_160;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h20 == lineSel) begin
            dirty_32 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_33 <= _GEN_161;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h21 == lineSel) begin
            dirty_33 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_34 <= _GEN_162;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h22 == lineSel) begin
            dirty_34 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_35 <= _GEN_163;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h23 == lineSel) begin
            dirty_35 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_36 <= _GEN_164;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h24 == lineSel) begin
            dirty_36 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_37 <= _GEN_165;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h25 == lineSel) begin
            dirty_37 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_38 <= _GEN_166;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h26 == lineSel) begin
            dirty_38 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_39 <= _GEN_167;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h27 == lineSel) begin
            dirty_39 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_40 <= _GEN_168;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h28 == lineSel) begin
            dirty_40 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_41 <= _GEN_169;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h29 == lineSel) begin
            dirty_41 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_42 <= _GEN_170;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h2a == lineSel) begin
            dirty_42 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_43 <= _GEN_171;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h2b == lineSel) begin
            dirty_43 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_44 <= _GEN_172;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h2c == lineSel) begin
            dirty_44 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_45 <= _GEN_173;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h2d == lineSel) begin
            dirty_45 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_46 <= _GEN_174;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h2e == lineSel) begin
            dirty_46 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_47 <= _GEN_175;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h2f == lineSel) begin
            dirty_47 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_48 <= _GEN_176;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h30 == lineSel) begin
            dirty_48 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_49 <= _GEN_177;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h31 == lineSel) begin
            dirty_49 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_50 <= _GEN_178;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h32 == lineSel) begin
            dirty_50 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_51 <= _GEN_179;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h33 == lineSel) begin
            dirty_51 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_52 <= _GEN_180;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h34 == lineSel) begin
            dirty_52 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_53 <= _GEN_181;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h35 == lineSel) begin
            dirty_53 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_54 <= _GEN_182;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h36 == lineSel) begin
            dirty_54 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_55 <= _GEN_183;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h37 == lineSel) begin
            dirty_55 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_56 <= _GEN_184;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h38 == lineSel) begin
            dirty_56 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_57 <= _GEN_185;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h39 == lineSel) begin
            dirty_57 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_58 <= _GEN_186;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h3a == lineSel) begin
            dirty_58 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_59 <= _GEN_187;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h3b == lineSel) begin
            dirty_59 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_60 <= _GEN_188;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h3c == lineSel) begin
            dirty_60 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_61 <= _GEN_189;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h3d == lineSel) begin
            dirty_61 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_62 <= _GEN_190;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h3e == lineSel) begin
            dirty_62 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_63 <= _GEN_191;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h3f == lineSel) begin
            dirty_63 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_64 <= _GEN_192;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h40 == lineSel) begin
            dirty_64 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_65 <= _GEN_193;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h41 == lineSel) begin
            dirty_65 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_66 <= _GEN_194;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h42 == lineSel) begin
            dirty_66 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_67 <= _GEN_195;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h43 == lineSel) begin
            dirty_67 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_68 <= _GEN_196;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h44 == lineSel) begin
            dirty_68 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_69 <= _GEN_197;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h45 == lineSel) begin
            dirty_69 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_70 <= _GEN_198;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h46 == lineSel) begin
            dirty_70 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_71 <= _GEN_199;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h47 == lineSel) begin
            dirty_71 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_72 <= _GEN_200;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h48 == lineSel) begin
            dirty_72 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_73 <= _GEN_201;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h49 == lineSel) begin
            dirty_73 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_74 <= _GEN_202;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h4a == lineSel) begin
            dirty_74 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_75 <= _GEN_203;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h4b == lineSel) begin
            dirty_75 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_76 <= _GEN_204;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h4c == lineSel) begin
            dirty_76 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_77 <= _GEN_205;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h4d == lineSel) begin
            dirty_77 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_78 <= _GEN_206;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h4e == lineSel) begin
            dirty_78 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_79 <= _GEN_207;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h4f == lineSel) begin
            dirty_79 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_80 <= _GEN_208;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h50 == lineSel) begin
            dirty_80 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_81 <= _GEN_209;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h51 == lineSel) begin
            dirty_81 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_82 <= _GEN_210;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h52 == lineSel) begin
            dirty_82 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_83 <= _GEN_211;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h53 == lineSel) begin
            dirty_83 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_84 <= _GEN_212;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h54 == lineSel) begin
            dirty_84 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_85 <= _GEN_213;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h55 == lineSel) begin
            dirty_85 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_86 <= _GEN_214;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h56 == lineSel) begin
            dirty_86 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_87 <= _GEN_215;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h57 == lineSel) begin
            dirty_87 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_88 <= _GEN_216;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h58 == lineSel) begin
            dirty_88 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_89 <= _GEN_217;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h59 == lineSel) begin
            dirty_89 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_90 <= _GEN_218;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h5a == lineSel) begin
            dirty_90 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_91 <= _GEN_219;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h5b == lineSel) begin
            dirty_91 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_92 <= _GEN_220;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h5c == lineSel) begin
            dirty_92 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_93 <= _GEN_221;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h5d == lineSel) begin
            dirty_93 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_94 <= _GEN_222;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h5e == lineSel) begin
            dirty_94 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_95 <= _GEN_223;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h5f == lineSel) begin
            dirty_95 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_96 <= _GEN_224;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h60 == lineSel) begin
            dirty_96 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_97 <= _GEN_225;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h61 == lineSel) begin
            dirty_97 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_98 <= _GEN_226;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h62 == lineSel) begin
            dirty_98 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_99 <= _GEN_227;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h63 == lineSel) begin
            dirty_99 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_100 <= _GEN_228;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h64 == lineSel) begin
            dirty_100 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_101 <= _GEN_229;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h65 == lineSel) begin
            dirty_101 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_102 <= _GEN_230;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h66 == lineSel) begin
            dirty_102 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_103 <= _GEN_231;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h67 == lineSel) begin
            dirty_103 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_104 <= _GEN_232;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h68 == lineSel) begin
            dirty_104 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_105 <= _GEN_233;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h69 == lineSel) begin
            dirty_105 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_106 <= _GEN_234;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h6a == lineSel) begin
            dirty_106 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_107 <= _GEN_235;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h6b == lineSel) begin
            dirty_107 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_108 <= _GEN_236;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h6c == lineSel) begin
            dirty_108 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_109 <= _GEN_237;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h6d == lineSel) begin
            dirty_109 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_110 <= _GEN_238;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h6e == lineSel) begin
            dirty_110 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_111 <= _GEN_239;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h6f == lineSel) begin
            dirty_111 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_112 <= _GEN_240;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h70 == lineSel) begin
            dirty_112 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_113 <= _GEN_241;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h71 == lineSel) begin
            dirty_113 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_114 <= _GEN_242;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h72 == lineSel) begin
            dirty_114 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_115 <= _GEN_243;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h73 == lineSel) begin
            dirty_115 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_116 <= _GEN_244;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h74 == lineSel) begin
            dirty_116 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_117 <= _GEN_245;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h75 == lineSel) begin
            dirty_117 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_118 <= _GEN_246;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h76 == lineSel) begin
            dirty_118 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_119 <= _GEN_247;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h77 == lineSel) begin
            dirty_119 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_120 <= _GEN_248;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h78 == lineSel) begin
            dirty_120 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_121 <= _GEN_249;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h79 == lineSel) begin
            dirty_121 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_122 <= _GEN_250;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h7a == lineSel) begin
            dirty_122 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_123 <= _GEN_251;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h7b == lineSel) begin
            dirty_123 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_124 <= _GEN_252;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h7c == lineSel) begin
            dirty_124 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_125 <= _GEN_253;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h7d == lineSel) begin
            dirty_125 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_126 <= _GEN_254;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h7e == lineSel) begin
            dirty_126 <= 1'h0;
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (cacheHit) begin
            if (_T_276) begin
              dirty_127 <= _GEN_255;
            end
          end
        end
      end
    end else if (!(_T_278)) begin
      if (_T_280) begin
        if (_T_283) begin
          if (7'h7f == lineSel) begin
            dirty_127 <= 1'h0;
          end
        end
      end
    end
    if (!(_T_274)) begin
      if (_T_278) begin
        if (_T_279) begin
          dataOffset <= 5'h0;
        end
      end else if (_T_280) begin
        if (io_axi_readData_valid) begin
          dataOffset <= _T_282;
        end
      end else if (!(_T_285)) begin
        if (_T_286) begin
          if (_T_287) begin
            dataOffset <= 5'h0;
          end
        end else if (_T_288) begin
          if (_T_290) begin
            dataOffset <= _T_282;
          end else begin
            dataOffset <= lastOffset;
          end
        end else if (_T_293) begin
          if (_T_287) begin
            dataOffset <= 5'h0;
          end
        end else if (_T_295) begin
          if (_T_290) begin
            dataOffset <= _T_282;
          end
        end
      end
    end
    if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (!(_T_280)) begin
          if (!(_T_285)) begin
            if (_T_286) begin
              if (_T_287) begin
                lastOffset <= 5'h0;
              end
            end else if (_T_288) begin
              if (_T_290) begin
                lastOffset <= dataOffset;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      aren <= 1'h0;
    end else if (!(_T_274)) begin
      if (_T_278) begin
        if (_T_279) begin
          aren <= 1'h0;
        end else begin
          aren <= 1'h1;
        end
      end
    end
    if (!(_T_274)) begin
      if (_T_278) begin
        raddr <= startRaddr;
      end
    end
    if (reset) begin
      awen <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (!(_T_280)) begin
          if (!(_T_285)) begin
            if (_T_286) begin
              if (_T_287) begin
                awen <= 1'h0;
              end else begin
                awen <= 1'h1;
              end
            end else if (!(_T_288)) begin
              if (_T_293) begin
                if (_T_287) begin
                  awen <= 1'h0;
                end else begin
                  awen <= 1'h1;
                end
              end
            end
          end
        end
      end
    end
    if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (!(_T_280)) begin
          if (!(_T_285)) begin
            if (_T_286) begin
              waddr <= startWaddr;
            end else if (!(_T_288)) begin
              if (_T_293) begin
                waddr <= flushAddr;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      wen <= 1'h0;
    end else if (!(_T_274)) begin
      if (!(_T_278)) begin
        if (!(_T_280)) begin
          if (!(_T_285)) begin
            if (!(_T_286)) begin
              if (_T_288) begin
                if (wlast) begin
                  wen <= 1'h0;
                end else begin
                  wen <= _T_290;
                end
              end else if (!(_T_293)) begin
                if (_T_295) begin
                  if (wlast) begin
                    wen <= 1'h0;
                  end else begin
                    wen <= _T_290;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_274) begin
      if (!(_T_275)) begin
        if (io_sram_en) begin
          if (!(cacheHit)) begin
            sramAddr <= io_sram_addr;
          end
        end
      end
    end
  end
endmodule
module Uncached(
  input         clock,
  input         reset,
  input         io_sram_en,
  output        io_sram_valid,
  input  [3:0]  io_sram_wen,
  input  [31:0] io_sram_addr,
  output [31:0] io_sram_rdata,
  input  [31:0] io_sram_wdata,
  input         io_axi_readAddr_ready,
  output        io_axi_readAddr_valid,
  output [31:0] io_axi_readAddr_bits_addr,
  input         io_axi_readData_valid,
  input  [31:0] io_axi_readData_bits_data,
  input         io_axi_readData_bits_last,
  input         io_axi_writeAddr_ready,
  output        io_axi_writeAddr_valid,
  output [31:0] io_axi_writeAddr_bits_addr,
  input         io_axi_writeData_ready,
  output        io_axi_writeData_valid,
  output [31:0] io_axi_writeData_bits_data,
  output        io_axi_writeData_bits_last,
  output [3:0]  io_axi_writeData_bits_strb
);
  reg [2:0] state; // @[Uncached.scala 25:22]
  reg [31:0] _RAND_0;
  reg [31:0] rdata; // @[Uncached.scala 28:20]
  reg [31:0] _RAND_1;
  wire  rvalid = io_axi_readData_valid & io_axi_readData_bits_last; // @[Uncached.scala 31:39]
  wire  _T = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_1 = io_sram_wen != 4'h0; // @[Uncached.scala 38:34]
  wire  _T_3 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_5 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_6 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_7 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_8 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_9 = state == 3'h6; // @[Uncached.scala 71:26]
  assign io_sram_valid = _T_9 | rvalid; // @[Uncached.scala 71:17]
  assign io_sram_rdata = rdata; // @[Uncached.scala 73:17]
  assign io_axi_readAddr_valid = state == 3'h1; // @[AXI.scala 56:20 Uncached.scala 77:31]
  assign io_axi_readAddr_bits_addr = io_sram_addr; // @[AXI.scala 9:21 Uncached.scala 78:31]
  assign io_axi_writeAddr_valid = state == 3'h3; // @[AXI.scala 59:21 Uncached.scala 82:31]
  assign io_axi_writeAddr_bits_addr = io_sram_addr; // @[AXI.scala 9:21 Uncached.scala 83:31]
  assign io_axi_writeData_valid = state == 3'h4; // @[AXI.scala 61:21 Uncached.scala 85:31]
  assign io_axi_writeData_bits_data = io_sram_wdata; // @[AXI.scala 9:21 Uncached.scala 86:31]
  assign io_axi_writeData_bits_last = state == 3'h4; // @[AXI.scala 9:21 Uncached.scala 87:31]
  assign io_axi_writeData_bits_strb = io_sram_wen; // @[AXI.scala 9:21 Uncached.scala 88:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  rdata = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (_T) begin
      if (io_sram_en) begin
        if (_T_1) begin
          state <= 3'h3;
        end else begin
          state <= 3'h1;
        end
      end
    end else if (_T_3) begin
      if (io_axi_readAddr_ready) begin
        state <= 3'h2;
      end
    end else if (_T_4) begin
      if (rvalid) begin
        state <= 3'h5;
      end
    end else if (_T_5) begin
      if (io_axi_writeAddr_ready) begin
        state <= 3'h4;
      end
    end else if (_T_6) begin
      if (io_axi_writeData_ready) begin
        state <= 3'h6;
      end
    end else if (_T_7) begin
      state <= 3'h0;
    end else if (_T_8) begin
      state <= 3'h0;
    end
    if (!(_T)) begin
      if (!(_T_3)) begin
        if (_T_4) begin
          if (rvalid) begin
            rdata <= io_axi_readData_bits_data;
          end
        end
      end
    end
  end
endmodule
module CoreBus(
  input         clock,
  input         reset,
  output        io_rom_valid,
  output        io_rom_fault,
  input  [31:0] io_rom_addr,
  output [31:0] io_rom_rdata,
  input         io_ram_en,
  output        io_ram_valid,
  output        io_ram_fault,
  input  [3:0]  io_ram_wen,
  input  [31:0] io_ram_addr,
  output [31:0] io_ram_rdata,
  input  [31:0] io_ram_wdata,
  input         io_tlb_en,
  input         io_tlb_flushInst,
  input         io_tlb_flushData,
  input  [21:0] io_tlb_basePpn,
  input         io_tlb_sum,
  input         io_tlb_smode,
  input         io_cache_flushInst,
  input         io_cache_flushData,
  input         io_inst_readAddr_ready,
  output        io_inst_readAddr_valid,
  output [31:0] io_inst_readAddr_bits_addr,
  input         io_inst_readData_valid,
  input  [31:0] io_inst_readData_bits_data,
  input         io_inst_readData_bits_last,
  input         io_data_readAddr_ready,
  output        io_data_readAddr_valid,
  output [31:0] io_data_readAddr_bits_addr,
  input         io_data_readData_valid,
  input  [31:0] io_data_readData_bits_data,
  input         io_data_readData_bits_last,
  input         io_data_writeAddr_ready,
  output        io_data_writeAddr_valid,
  output [31:0] io_data_writeAddr_bits_addr,
  input         io_data_writeData_ready,
  output        io_data_writeData_valid,
  output [31:0] io_data_writeData_bits_data,
  output        io_data_writeData_bits_last,
  input         io_uncached_readAddr_ready,
  output        io_uncached_readAddr_valid,
  output [31:0] io_uncached_readAddr_bits_addr,
  input         io_uncached_readData_valid,
  input  [31:0] io_uncached_readData_bits_data,
  input         io_uncached_readData_bits_last,
  input         io_uncached_writeAddr_ready,
  output        io_uncached_writeAddr_valid,
  output [31:0] io_uncached_writeAddr_bits_addr,
  input         io_uncached_writeData_ready,
  output        io_uncached_writeData_valid,
  output [31:0] io_uncached_writeData_bits_data,
  output        io_uncached_writeData_bits_last,
  output [3:0]  io_uncached_writeData_bits_strb
);
  wire  immu_clock; // @[CoreBus.scala 64:20]
  wire  immu_reset; // @[CoreBus.scala 64:20]
  wire  immu_io_en; // @[CoreBus.scala 64:20]
  wire  immu_io_flush; // @[CoreBus.scala 64:20]
  wire [21:0] immu_io_basePpn; // @[CoreBus.scala 64:20]
  wire  immu_io_sum; // @[CoreBus.scala 64:20]
  wire  immu_io_smode; // @[CoreBus.scala 64:20]
  wire [31:0] immu_io_vaddr; // @[CoreBus.scala 64:20]
  wire  immu_io_valid; // @[CoreBus.scala 64:20]
  wire  immu_io_fault; // @[CoreBus.scala 64:20]
  wire [31:0] immu_io_paddr; // @[CoreBus.scala 64:20]
  wire  immu_io_data_en; // @[CoreBus.scala 64:20]
  wire  immu_io_data_valid; // @[CoreBus.scala 64:20]
  wire [31:0] immu_io_data_addr; // @[CoreBus.scala 64:20]
  wire [31:0] immu_io_data_rdata; // @[CoreBus.scala 64:20]
  wire  idemux_io_sel2; // @[CoreBus.scala 75:22]
  wire  idemux_io_in1_en; // @[CoreBus.scala 75:22]
  wire  idemux_io_in1_valid; // @[CoreBus.scala 75:22]
  wire [31:0] idemux_io_in1_addr; // @[CoreBus.scala 75:22]
  wire [31:0] idemux_io_in1_rdata; // @[CoreBus.scala 75:22]
  wire  idemux_io_in2_en; // @[CoreBus.scala 75:22]
  wire  idemux_io_in2_valid; // @[CoreBus.scala 75:22]
  wire [3:0] idemux_io_in2_wen; // @[CoreBus.scala 75:22]
  wire [31:0] idemux_io_in2_addr; // @[CoreBus.scala 75:22]
  wire [31:0] idemux_io_in2_rdata; // @[CoreBus.scala 75:22]
  wire [31:0] idemux_io_in2_wdata; // @[CoreBus.scala 75:22]
  wire  idemux_io_out_en; // @[CoreBus.scala 75:22]
  wire  idemux_io_out_valid; // @[CoreBus.scala 75:22]
  wire [3:0] idemux_io_out_wen; // @[CoreBus.scala 75:22]
  wire [31:0] idemux_io_out_addr; // @[CoreBus.scala 75:22]
  wire [31:0] idemux_io_out_rdata; // @[CoreBus.scala 75:22]
  wire [31:0] idemux_io_out_wdata; // @[CoreBus.scala 75:22]
  wire  icache_clock; // @[CoreBus.scala 82:22]
  wire  icache_reset; // @[CoreBus.scala 82:22]
  wire  icache_io_sram_en; // @[CoreBus.scala 82:22]
  wire  icache_io_sram_valid; // @[CoreBus.scala 82:22]
  wire [31:0] icache_io_sram_addr; // @[CoreBus.scala 82:22]
  wire [31:0] icache_io_sram_rdata; // @[CoreBus.scala 82:22]
  wire  icache_io_flush; // @[CoreBus.scala 82:22]
  wire  icache_io_axi_readAddr_ready; // @[CoreBus.scala 82:22]
  wire  icache_io_axi_readAddr_valid; // @[CoreBus.scala 82:22]
  wire [31:0] icache_io_axi_readAddr_bits_addr; // @[CoreBus.scala 82:22]
  wire  icache_io_axi_readData_valid; // @[CoreBus.scala 82:22]
  wire [31:0] icache_io_axi_readData_bits_data; // @[CoreBus.scala 82:22]
  wire  icache_io_axi_readData_bits_last; // @[CoreBus.scala 82:22]
  wire  dmmu_clock; // @[CoreBus.scala 91:20]
  wire  dmmu_reset; // @[CoreBus.scala 91:20]
  wire  dmmu_io_en; // @[CoreBus.scala 91:20]
  wire  dmmu_io_flush; // @[CoreBus.scala 91:20]
  wire [21:0] dmmu_io_basePpn; // @[CoreBus.scala 91:20]
  wire  dmmu_io_sum; // @[CoreBus.scala 91:20]
  wire  dmmu_io_smode; // @[CoreBus.scala 91:20]
  wire  dmmu_io_lookup; // @[CoreBus.scala 91:20]
  wire  dmmu_io_write; // @[CoreBus.scala 91:20]
  wire [31:0] dmmu_io_vaddr; // @[CoreBus.scala 91:20]
  wire  dmmu_io_valid; // @[CoreBus.scala 91:20]
  wire  dmmu_io_fault; // @[CoreBus.scala 91:20]
  wire [31:0] dmmu_io_paddr; // @[CoreBus.scala 91:20]
  wire  dmmu_io_data_en; // @[CoreBus.scala 91:20]
  wire  dmmu_io_data_valid; // @[CoreBus.scala 91:20]
  wire [31:0] dmmu_io_data_addr; // @[CoreBus.scala 91:20]
  wire [31:0] dmmu_io_data_rdata; // @[CoreBus.scala 91:20]
  wire  ddemux_io_sel2; // @[CoreBus.scala 102:22]
  wire  ddemux_io_in1_en; // @[CoreBus.scala 102:22]
  wire  ddemux_io_in1_valid; // @[CoreBus.scala 102:22]
  wire [31:0] ddemux_io_in1_addr; // @[CoreBus.scala 102:22]
  wire [31:0] ddemux_io_in1_rdata; // @[CoreBus.scala 102:22]
  wire  ddemux_io_in2_en; // @[CoreBus.scala 102:22]
  wire  ddemux_io_in2_valid; // @[CoreBus.scala 102:22]
  wire [3:0] ddemux_io_in2_wen; // @[CoreBus.scala 102:22]
  wire [31:0] ddemux_io_in2_addr; // @[CoreBus.scala 102:22]
  wire [31:0] ddemux_io_in2_rdata; // @[CoreBus.scala 102:22]
  wire [31:0] ddemux_io_in2_wdata; // @[CoreBus.scala 102:22]
  wire  ddemux_io_out_en; // @[CoreBus.scala 102:22]
  wire  ddemux_io_out_valid; // @[CoreBus.scala 102:22]
  wire [3:0] ddemux_io_out_wen; // @[CoreBus.scala 102:22]
  wire [31:0] ddemux_io_out_addr; // @[CoreBus.scala 102:22]
  wire [31:0] ddemux_io_out_rdata; // @[CoreBus.scala 102:22]
  wire [31:0] ddemux_io_out_wdata; // @[CoreBus.scala 102:22]
  wire  mux_clock; // @[CoreBus.scala 109:19]
  wire  mux_io_sel2; // @[CoreBus.scala 109:19]
  wire  mux_io_in_en; // @[CoreBus.scala 109:19]
  wire  mux_io_in_valid; // @[CoreBus.scala 109:19]
  wire [3:0] mux_io_in_wen; // @[CoreBus.scala 109:19]
  wire [31:0] mux_io_in_addr; // @[CoreBus.scala 109:19]
  wire [31:0] mux_io_in_rdata; // @[CoreBus.scala 109:19]
  wire [31:0] mux_io_in_wdata; // @[CoreBus.scala 109:19]
  wire  mux_io_out1_en; // @[CoreBus.scala 109:19]
  wire  mux_io_out1_valid; // @[CoreBus.scala 109:19]
  wire [3:0] mux_io_out1_wen; // @[CoreBus.scala 109:19]
  wire [31:0] mux_io_out1_addr; // @[CoreBus.scala 109:19]
  wire [31:0] mux_io_out1_rdata; // @[CoreBus.scala 109:19]
  wire [31:0] mux_io_out1_wdata; // @[CoreBus.scala 109:19]
  wire  mux_io_out2_en; // @[CoreBus.scala 109:19]
  wire  mux_io_out2_valid; // @[CoreBus.scala 109:19]
  wire [3:0] mux_io_out2_wen; // @[CoreBus.scala 109:19]
  wire [31:0] mux_io_out2_addr; // @[CoreBus.scala 109:19]
  wire [31:0] mux_io_out2_rdata; // @[CoreBus.scala 109:19]
  wire [31:0] mux_io_out2_wdata; // @[CoreBus.scala 109:19]
  wire  dcache_clock; // @[CoreBus.scala 115:22]
  wire  dcache_reset; // @[CoreBus.scala 115:22]
  wire  dcache_io_sram_en; // @[CoreBus.scala 115:22]
  wire  dcache_io_sram_valid; // @[CoreBus.scala 115:22]
  wire [3:0] dcache_io_sram_wen; // @[CoreBus.scala 115:22]
  wire [31:0] dcache_io_sram_addr; // @[CoreBus.scala 115:22]
  wire [31:0] dcache_io_sram_rdata; // @[CoreBus.scala 115:22]
  wire [31:0] dcache_io_sram_wdata; // @[CoreBus.scala 115:22]
  wire  dcache_io_flush; // @[CoreBus.scala 115:22]
  wire  dcache_io_axi_readAddr_ready; // @[CoreBus.scala 115:22]
  wire  dcache_io_axi_readAddr_valid; // @[CoreBus.scala 115:22]
  wire [31:0] dcache_io_axi_readAddr_bits_addr; // @[CoreBus.scala 115:22]
  wire  dcache_io_axi_readData_valid; // @[CoreBus.scala 115:22]
  wire [31:0] dcache_io_axi_readData_bits_data; // @[CoreBus.scala 115:22]
  wire  dcache_io_axi_readData_bits_last; // @[CoreBus.scala 115:22]
  wire  dcache_io_axi_writeAddr_ready; // @[CoreBus.scala 115:22]
  wire  dcache_io_axi_writeAddr_valid; // @[CoreBus.scala 115:22]
  wire [31:0] dcache_io_axi_writeAddr_bits_addr; // @[CoreBus.scala 115:22]
  wire  dcache_io_axi_writeData_ready; // @[CoreBus.scala 115:22]
  wire  dcache_io_axi_writeData_valid; // @[CoreBus.scala 115:22]
  wire [31:0] dcache_io_axi_writeData_bits_data; // @[CoreBus.scala 115:22]
  wire  dcache_io_axi_writeData_bits_last; // @[CoreBus.scala 115:22]
  wire  uncached_clock; // @[CoreBus.scala 121:24]
  wire  uncached_reset; // @[CoreBus.scala 121:24]
  wire  uncached_io_sram_en; // @[CoreBus.scala 121:24]
  wire  uncached_io_sram_valid; // @[CoreBus.scala 121:24]
  wire [3:0] uncached_io_sram_wen; // @[CoreBus.scala 121:24]
  wire [31:0] uncached_io_sram_addr; // @[CoreBus.scala 121:24]
  wire [31:0] uncached_io_sram_rdata; // @[CoreBus.scala 121:24]
  wire [31:0] uncached_io_sram_wdata; // @[CoreBus.scala 121:24]
  wire  uncached_io_axi_readAddr_ready; // @[CoreBus.scala 121:24]
  wire  uncached_io_axi_readAddr_valid; // @[CoreBus.scala 121:24]
  wire [31:0] uncached_io_axi_readAddr_bits_addr; // @[CoreBus.scala 121:24]
  wire  uncached_io_axi_readData_valid; // @[CoreBus.scala 121:24]
  wire [31:0] uncached_io_axi_readData_bits_data; // @[CoreBus.scala 121:24]
  wire  uncached_io_axi_readData_bits_last; // @[CoreBus.scala 121:24]
  wire  uncached_io_axi_writeAddr_ready; // @[CoreBus.scala 121:24]
  wire  uncached_io_axi_writeAddr_valid; // @[CoreBus.scala 121:24]
  wire [31:0] uncached_io_axi_writeAddr_bits_addr; // @[CoreBus.scala 121:24]
  wire  uncached_io_axi_writeData_ready; // @[CoreBus.scala 121:24]
  wire  uncached_io_axi_writeData_valid; // @[CoreBus.scala 121:24]
  wire [31:0] uncached_io_axi_writeData_bits_data; // @[CoreBus.scala 121:24]
  wire  uncached_io_axi_writeData_bits_last; // @[CoreBus.scala 121:24]
  wire [3:0] uncached_io_axi_writeData_bits_strb; // @[CoreBus.scala 121:24]
  wire  _T_2 = dmmu_io_paddr >= 32'h10000000; // @[CoreBus.scala 110:32]
  wire  _T_3 = dmmu_io_paddr < 32'h20000000; // @[CoreBus.scala 111:32]
  MMU immu ( // @[CoreBus.scala 64:20]
    .clock(immu_clock),
    .reset(immu_reset),
    .io_en(immu_io_en),
    .io_flush(immu_io_flush),
    .io_basePpn(immu_io_basePpn),
    .io_sum(immu_io_sum),
    .io_smode(immu_io_smode),
    .io_vaddr(immu_io_vaddr),
    .io_valid(immu_io_valid),
    .io_fault(immu_io_fault),
    .io_paddr(immu_io_paddr),
    .io_data_en(immu_io_data_en),
    .io_data_valid(immu_io_data_valid),
    .io_data_addr(immu_io_data_addr),
    .io_data_rdata(immu_io_data_rdata)
  );
  SramDemux2 idemux ( // @[CoreBus.scala 75:22]
    .io_sel2(idemux_io_sel2),
    .io_in1_en(idemux_io_in1_en),
    .io_in1_valid(idemux_io_in1_valid),
    .io_in1_addr(idemux_io_in1_addr),
    .io_in1_rdata(idemux_io_in1_rdata),
    .io_in2_en(idemux_io_in2_en),
    .io_in2_valid(idemux_io_in2_valid),
    .io_in2_wen(idemux_io_in2_wen),
    .io_in2_addr(idemux_io_in2_addr),
    .io_in2_rdata(idemux_io_in2_rdata),
    .io_in2_wdata(idemux_io_in2_wdata),
    .io_out_en(idemux_io_out_en),
    .io_out_valid(idemux_io_out_valid),
    .io_out_wen(idemux_io_out_wen),
    .io_out_addr(idemux_io_out_addr),
    .io_out_rdata(idemux_io_out_rdata),
    .io_out_wdata(idemux_io_out_wdata)
  );
  InstCache icache ( // @[CoreBus.scala 82:22]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_sram_en(icache_io_sram_en),
    .io_sram_valid(icache_io_sram_valid),
    .io_sram_addr(icache_io_sram_addr),
    .io_sram_rdata(icache_io_sram_rdata),
    .io_flush(icache_io_flush),
    .io_axi_readAddr_ready(icache_io_axi_readAddr_ready),
    .io_axi_readAddr_valid(icache_io_axi_readAddr_valid),
    .io_axi_readAddr_bits_addr(icache_io_axi_readAddr_bits_addr),
    .io_axi_readData_valid(icache_io_axi_readData_valid),
    .io_axi_readData_bits_data(icache_io_axi_readData_bits_data),
    .io_axi_readData_bits_last(icache_io_axi_readData_bits_last)
  );
  MMU_1 dmmu ( // @[CoreBus.scala 91:20]
    .clock(dmmu_clock),
    .reset(dmmu_reset),
    .io_en(dmmu_io_en),
    .io_flush(dmmu_io_flush),
    .io_basePpn(dmmu_io_basePpn),
    .io_sum(dmmu_io_sum),
    .io_smode(dmmu_io_smode),
    .io_lookup(dmmu_io_lookup),
    .io_write(dmmu_io_write),
    .io_vaddr(dmmu_io_vaddr),
    .io_valid(dmmu_io_valid),
    .io_fault(dmmu_io_fault),
    .io_paddr(dmmu_io_paddr),
    .io_data_en(dmmu_io_data_en),
    .io_data_valid(dmmu_io_data_valid),
    .io_data_addr(dmmu_io_data_addr),
    .io_data_rdata(dmmu_io_data_rdata)
  );
  SramDemux2 ddemux ( // @[CoreBus.scala 102:22]
    .io_sel2(ddemux_io_sel2),
    .io_in1_en(ddemux_io_in1_en),
    .io_in1_valid(ddemux_io_in1_valid),
    .io_in1_addr(ddemux_io_in1_addr),
    .io_in1_rdata(ddemux_io_in1_rdata),
    .io_in2_en(ddemux_io_in2_en),
    .io_in2_valid(ddemux_io_in2_valid),
    .io_in2_wen(ddemux_io_in2_wen),
    .io_in2_addr(ddemux_io_in2_addr),
    .io_in2_rdata(ddemux_io_in2_rdata),
    .io_in2_wdata(ddemux_io_in2_wdata),
    .io_out_en(ddemux_io_out_en),
    .io_out_valid(ddemux_io_out_valid),
    .io_out_wen(ddemux_io_out_wen),
    .io_out_addr(ddemux_io_out_addr),
    .io_out_rdata(ddemux_io_out_rdata),
    .io_out_wdata(ddemux_io_out_wdata)
  );
  SramMux2 mux ( // @[CoreBus.scala 109:19]
    .clock(mux_clock),
    .io_sel2(mux_io_sel2),
    .io_in_en(mux_io_in_en),
    .io_in_valid(mux_io_in_valid),
    .io_in_wen(mux_io_in_wen),
    .io_in_addr(mux_io_in_addr),
    .io_in_rdata(mux_io_in_rdata),
    .io_in_wdata(mux_io_in_wdata),
    .io_out1_en(mux_io_out1_en),
    .io_out1_valid(mux_io_out1_valid),
    .io_out1_wen(mux_io_out1_wen),
    .io_out1_addr(mux_io_out1_addr),
    .io_out1_rdata(mux_io_out1_rdata),
    .io_out1_wdata(mux_io_out1_wdata),
    .io_out2_en(mux_io_out2_en),
    .io_out2_valid(mux_io_out2_valid),
    .io_out2_wen(mux_io_out2_wen),
    .io_out2_addr(mux_io_out2_addr),
    .io_out2_rdata(mux_io_out2_rdata),
    .io_out2_wdata(mux_io_out2_wdata)
  );
  DataCache dcache ( // @[CoreBus.scala 115:22]
    .clock(dcache_clock),
    .reset(dcache_reset),
    .io_sram_en(dcache_io_sram_en),
    .io_sram_valid(dcache_io_sram_valid),
    .io_sram_wen(dcache_io_sram_wen),
    .io_sram_addr(dcache_io_sram_addr),
    .io_sram_rdata(dcache_io_sram_rdata),
    .io_sram_wdata(dcache_io_sram_wdata),
    .io_flush(dcache_io_flush),
    .io_axi_readAddr_ready(dcache_io_axi_readAddr_ready),
    .io_axi_readAddr_valid(dcache_io_axi_readAddr_valid),
    .io_axi_readAddr_bits_addr(dcache_io_axi_readAddr_bits_addr),
    .io_axi_readData_valid(dcache_io_axi_readData_valid),
    .io_axi_readData_bits_data(dcache_io_axi_readData_bits_data),
    .io_axi_readData_bits_last(dcache_io_axi_readData_bits_last),
    .io_axi_writeAddr_ready(dcache_io_axi_writeAddr_ready),
    .io_axi_writeAddr_valid(dcache_io_axi_writeAddr_valid),
    .io_axi_writeAddr_bits_addr(dcache_io_axi_writeAddr_bits_addr),
    .io_axi_writeData_ready(dcache_io_axi_writeData_ready),
    .io_axi_writeData_valid(dcache_io_axi_writeData_valid),
    .io_axi_writeData_bits_data(dcache_io_axi_writeData_bits_data),
    .io_axi_writeData_bits_last(dcache_io_axi_writeData_bits_last)
  );
  Uncached uncached ( // @[CoreBus.scala 121:24]
    .clock(uncached_clock),
    .reset(uncached_reset),
    .io_sram_en(uncached_io_sram_en),
    .io_sram_valid(uncached_io_sram_valid),
    .io_sram_wen(uncached_io_sram_wen),
    .io_sram_addr(uncached_io_sram_addr),
    .io_sram_rdata(uncached_io_sram_rdata),
    .io_sram_wdata(uncached_io_sram_wdata),
    .io_axi_readAddr_ready(uncached_io_axi_readAddr_ready),
    .io_axi_readAddr_valid(uncached_io_axi_readAddr_valid),
    .io_axi_readAddr_bits_addr(uncached_io_axi_readAddr_bits_addr),
    .io_axi_readData_valid(uncached_io_axi_readData_valid),
    .io_axi_readData_bits_data(uncached_io_axi_readData_bits_data),
    .io_axi_readData_bits_last(uncached_io_axi_readData_bits_last),
    .io_axi_writeAddr_ready(uncached_io_axi_writeAddr_ready),
    .io_axi_writeAddr_valid(uncached_io_axi_writeAddr_valid),
    .io_axi_writeAddr_bits_addr(uncached_io_axi_writeAddr_bits_addr),
    .io_axi_writeData_ready(uncached_io_axi_writeData_ready),
    .io_axi_writeData_valid(uncached_io_axi_writeData_valid),
    .io_axi_writeData_bits_data(uncached_io_axi_writeData_bits_data),
    .io_axi_writeData_bits_last(uncached_io_axi_writeData_bits_last),
    .io_axi_writeData_bits_strb(uncached_io_axi_writeData_bits_strb)
  );
  assign io_rom_valid = idemux_io_in2_valid; // @[CoreBus.scala 78:23]
  assign io_rom_fault = immu_io_fault; // @[CoreBus.scala 78:23 CoreBus.scala 88:17]
  assign io_rom_rdata = idemux_io_in2_rdata; // @[CoreBus.scala 78:23]
  assign io_ram_valid = ddemux_io_in2_valid; // @[CoreBus.scala 105:23]
  assign io_ram_fault = dmmu_io_fault; // @[CoreBus.scala 105:23 CoreBus.scala 126:17]
  assign io_ram_rdata = ddemux_io_in2_rdata; // @[CoreBus.scala 105:23]
  assign io_inst_readAddr_valid = icache_io_axi_readAddr_valid; // @[CoreBus.scala 85:19]
  assign io_inst_readAddr_bits_addr = icache_io_axi_readAddr_bits_addr; // @[CoreBus.scala 85:19]
  assign io_data_readAddr_valid = dcache_io_axi_readAddr_valid; // @[CoreBus.scala 118:19]
  assign io_data_readAddr_bits_addr = dcache_io_axi_readAddr_bits_addr; // @[CoreBus.scala 118:19]
  assign io_data_writeAddr_valid = dcache_io_axi_writeAddr_valid; // @[CoreBus.scala 118:19]
  assign io_data_writeAddr_bits_addr = dcache_io_axi_writeAddr_bits_addr; // @[CoreBus.scala 118:19]
  assign io_data_writeData_valid = dcache_io_axi_writeData_valid; // @[CoreBus.scala 118:19]
  assign io_data_writeData_bits_data = dcache_io_axi_writeData_bits_data; // @[CoreBus.scala 118:19]
  assign io_data_writeData_bits_last = dcache_io_axi_writeData_bits_last; // @[CoreBus.scala 118:19]
  assign io_uncached_readAddr_valid = uncached_io_axi_readAddr_valid; // @[CoreBus.scala 123:21]
  assign io_uncached_readAddr_bits_addr = uncached_io_axi_readAddr_bits_addr; // @[CoreBus.scala 123:21]
  assign io_uncached_writeAddr_valid = uncached_io_axi_writeAddr_valid; // @[CoreBus.scala 123:21]
  assign io_uncached_writeAddr_bits_addr = uncached_io_axi_writeAddr_bits_addr; // @[CoreBus.scala 123:21]
  assign io_uncached_writeData_valid = uncached_io_axi_writeData_valid; // @[CoreBus.scala 123:21]
  assign io_uncached_writeData_bits_data = uncached_io_axi_writeData_bits_data; // @[CoreBus.scala 123:21]
  assign io_uncached_writeData_bits_last = uncached_io_axi_writeData_bits_last; // @[CoreBus.scala 123:21]
  assign io_uncached_writeData_bits_strb = uncached_io_axi_writeData_bits_strb; // @[CoreBus.scala 123:21]
  assign immu_clock = clock;
  assign immu_reset = reset;
  assign immu_io_en = io_tlb_en; // @[CoreBus.scala 65:19]
  assign immu_io_flush = io_tlb_flushInst; // @[CoreBus.scala 66:19]
  assign immu_io_basePpn = io_tlb_basePpn; // @[CoreBus.scala 67:19]
  assign immu_io_sum = io_tlb_sum; // @[CoreBus.scala 68:19]
  assign immu_io_smode = io_tlb_smode; // @[CoreBus.scala 69:19]
  assign immu_io_vaddr = io_rom_addr; // @[CoreBus.scala 72:19]
  assign immu_io_data_valid = idemux_io_in1_valid; // @[CoreBus.scala 77:23]
  assign immu_io_data_rdata = idemux_io_in1_rdata; // @[CoreBus.scala 77:23]
  assign idemux_io_sel2 = immu_io_valid; // @[CoreBus.scala 76:23]
  assign idemux_io_in1_en = immu_io_data_en; // @[CoreBus.scala 77:23]
  assign idemux_io_in1_addr = immu_io_data_addr; // @[CoreBus.scala 77:23]
  assign idemux_io_in2_en = 1'h1; // @[CoreBus.scala 78:23]
  assign idemux_io_in2_wen = 4'h0; // @[CoreBus.scala 78:23]
  assign idemux_io_in2_addr = immu_io_paddr; // @[CoreBus.scala 78:23 CoreBus.scala 79:23]
  assign idemux_io_in2_wdata = 32'h0; // @[CoreBus.scala 78:23]
  assign idemux_io_out_valid = icache_io_sram_valid; // @[CoreBus.scala 83:19]
  assign idemux_io_out_rdata = icache_io_sram_rdata; // @[CoreBus.scala 83:19]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_sram_en = idemux_io_out_en; // @[CoreBus.scala 83:19]
  assign icache_io_sram_addr = idemux_io_out_addr; // @[CoreBus.scala 83:19]
  assign icache_io_flush = io_cache_flushInst; // @[CoreBus.scala 84:19]
  assign icache_io_axi_readAddr_ready = io_inst_readAddr_ready; // @[CoreBus.scala 85:19]
  assign icache_io_axi_readData_valid = io_inst_readData_valid; // @[CoreBus.scala 85:19]
  assign icache_io_axi_readData_bits_data = io_inst_readData_bits_data; // @[CoreBus.scala 85:19]
  assign icache_io_axi_readData_bits_last = io_inst_readData_bits_last; // @[CoreBus.scala 85:19]
  assign dmmu_clock = clock;
  assign dmmu_reset = reset;
  assign dmmu_io_en = io_tlb_en; // @[CoreBus.scala 92:19]
  assign dmmu_io_flush = io_tlb_flushData; // @[CoreBus.scala 93:19]
  assign dmmu_io_basePpn = io_tlb_basePpn; // @[CoreBus.scala 94:19]
  assign dmmu_io_sum = io_tlb_sum; // @[CoreBus.scala 95:19]
  assign dmmu_io_smode = io_tlb_smode; // @[CoreBus.scala 96:19]
  assign dmmu_io_lookup = io_ram_en; // @[CoreBus.scala 97:19]
  assign dmmu_io_write = io_ram_wen != 4'h0; // @[CoreBus.scala 98:19]
  assign dmmu_io_vaddr = io_ram_addr; // @[CoreBus.scala 99:19]
  assign dmmu_io_data_valid = ddemux_io_in1_valid; // @[CoreBus.scala 104:23]
  assign dmmu_io_data_rdata = ddemux_io_in1_rdata; // @[CoreBus.scala 104:23]
  assign ddemux_io_sel2 = dmmu_io_valid; // @[CoreBus.scala 103:23]
  assign ddemux_io_in1_en = dmmu_io_data_en; // @[CoreBus.scala 104:23]
  assign ddemux_io_in1_addr = dmmu_io_data_addr; // @[CoreBus.scala 104:23]
  assign ddemux_io_in2_en = io_ram_en; // @[CoreBus.scala 105:23]
  assign ddemux_io_in2_wen = io_ram_wen; // @[CoreBus.scala 105:23]
  assign ddemux_io_in2_addr = dmmu_io_paddr; // @[CoreBus.scala 105:23 CoreBus.scala 106:23]
  assign ddemux_io_in2_wdata = io_ram_wdata; // @[CoreBus.scala 105:23]
  assign ddemux_io_out_valid = mux_io_in_valid; // @[CoreBus.scala 112:15]
  assign ddemux_io_out_rdata = mux_io_in_rdata; // @[CoreBus.scala 112:15]
  assign mux_clock = clock;
  assign mux_io_sel2 = _T_2 & _T_3; // @[CoreBus.scala 110:15]
  assign mux_io_in_en = ddemux_io_out_en; // @[CoreBus.scala 112:15]
  assign mux_io_in_wen = ddemux_io_out_wen; // @[CoreBus.scala 112:15]
  assign mux_io_in_addr = ddemux_io_out_addr; // @[CoreBus.scala 112:15]
  assign mux_io_in_wdata = ddemux_io_out_wdata; // @[CoreBus.scala 112:15]
  assign mux_io_out1_valid = dcache_io_sram_valid; // @[CoreBus.scala 116:19]
  assign mux_io_out1_rdata = dcache_io_sram_rdata; // @[CoreBus.scala 116:19]
  assign mux_io_out2_valid = uncached_io_sram_valid; // @[CoreBus.scala 122:21]
  assign mux_io_out2_rdata = uncached_io_sram_rdata; // @[CoreBus.scala 122:21]
  assign dcache_clock = clock;
  assign dcache_reset = reset;
  assign dcache_io_sram_en = mux_io_out1_en; // @[CoreBus.scala 116:19]
  assign dcache_io_sram_wen = mux_io_out1_wen; // @[CoreBus.scala 116:19]
  assign dcache_io_sram_addr = mux_io_out1_addr; // @[CoreBus.scala 116:19]
  assign dcache_io_sram_wdata = mux_io_out1_wdata; // @[CoreBus.scala 116:19]
  assign dcache_io_flush = io_cache_flushData; // @[CoreBus.scala 117:19]
  assign dcache_io_axi_readAddr_ready = io_data_readAddr_ready; // @[CoreBus.scala 118:19]
  assign dcache_io_axi_readData_valid = io_data_readData_valid; // @[CoreBus.scala 118:19]
  assign dcache_io_axi_readData_bits_data = io_data_readData_bits_data; // @[CoreBus.scala 118:19]
  assign dcache_io_axi_readData_bits_last = io_data_readData_bits_last; // @[CoreBus.scala 118:19]
  assign dcache_io_axi_writeAddr_ready = io_data_writeAddr_ready; // @[CoreBus.scala 118:19]
  assign dcache_io_axi_writeData_ready = io_data_writeData_ready; // @[CoreBus.scala 118:19]
  assign uncached_clock = clock;
  assign uncached_reset = reset;
  assign uncached_io_sram_en = mux_io_out2_en; // @[CoreBus.scala 122:21]
  assign uncached_io_sram_wen = mux_io_out2_wen; // @[CoreBus.scala 122:21]
  assign uncached_io_sram_addr = mux_io_out2_addr; // @[CoreBus.scala 122:21]
  assign uncached_io_sram_wdata = mux_io_out2_wdata; // @[CoreBus.scala 122:21]
  assign uncached_io_axi_readAddr_ready = io_uncached_readAddr_ready; // @[CoreBus.scala 123:21]
  assign uncached_io_axi_readData_valid = io_uncached_readData_valid; // @[CoreBus.scala 123:21]
  assign uncached_io_axi_readData_bits_data = io_uncached_readData_bits_data; // @[CoreBus.scala 123:21]
  assign uncached_io_axi_readData_bits_last = io_uncached_readData_bits_last; // @[CoreBus.scala 123:21]
  assign uncached_io_axi_writeAddr_ready = io_uncached_writeAddr_ready; // @[CoreBus.scala 123:21]
  assign uncached_io_axi_writeData_ready = io_uncached_writeData_ready; // @[CoreBus.scala 123:21]
endmodule
module Fuxi(
  input         clock,
  input         reset,
  input         io_irq_timer,
  input         io_irq_soft,
  input         io_irq_extern,
  output        io_debug_regWen,
  output [4:0]  io_debug_regWaddr,
  output [31:0] io_debug_regWdata,
  output [31:0] io_debug_pc,
  input         io_inst_readAddr_ready,
  output        io_inst_readAddr_valid,
  output [31:0] io_inst_readAddr_bits_addr,
  output [3:0]  io_inst_readAddr_bits_id,
  output [2:0]  io_inst_readAddr_bits_size,
  output [7:0]  io_inst_readAddr_bits_len,
  output [1:0]  io_inst_readAddr_bits_burst,
  output        io_inst_readAddr_bits_lock,
  output [3:0]  io_inst_readAddr_bits_cache,
  output [2:0]  io_inst_readAddr_bits_prot,
  output        io_inst_readData_ready,
  input         io_inst_readData_valid,
  input  [31:0] io_inst_readData_bits_data,
  input  [3:0]  io_inst_readData_bits_id,
  input         io_inst_readData_bits_last,
  input  [1:0]  io_inst_readData_bits_resp,
  input         io_inst_writeAddr_ready,
  output        io_inst_writeAddr_valid,
  output [31:0] io_inst_writeAddr_bits_addr,
  output [3:0]  io_inst_writeAddr_bits_id,
  output [2:0]  io_inst_writeAddr_bits_size,
  output [7:0]  io_inst_writeAddr_bits_len,
  output [1:0]  io_inst_writeAddr_bits_burst,
  output        io_inst_writeAddr_bits_lock,
  output [3:0]  io_inst_writeAddr_bits_cache,
  output [2:0]  io_inst_writeAddr_bits_prot,
  input         io_inst_writeData_ready,
  output        io_inst_writeData_valid,
  output [31:0] io_inst_writeData_bits_data,
  output [3:0]  io_inst_writeData_bits_id,
  output        io_inst_writeData_bits_last,
  output [3:0]  io_inst_writeData_bits_strb,
  output        io_inst_writeResp_ready,
  input         io_inst_writeResp_valid,
  input  [3:0]  io_inst_writeResp_bits_id,
  input  [1:0]  io_inst_writeResp_bits_resp,
  input         io_data_readAddr_ready,
  output        io_data_readAddr_valid,
  output [31:0] io_data_readAddr_bits_addr,
  output [3:0]  io_data_readAddr_bits_id,
  output [2:0]  io_data_readAddr_bits_size,
  output [7:0]  io_data_readAddr_bits_len,
  output [1:0]  io_data_readAddr_bits_burst,
  output        io_data_readAddr_bits_lock,
  output [3:0]  io_data_readAddr_bits_cache,
  output [2:0]  io_data_readAddr_bits_prot,
  output        io_data_readData_ready,
  input         io_data_readData_valid,
  input  [31:0] io_data_readData_bits_data,
  input  [3:0]  io_data_readData_bits_id,
  input         io_data_readData_bits_last,
  input  [1:0]  io_data_readData_bits_resp,
  input         io_data_writeAddr_ready,
  output        io_data_writeAddr_valid,
  output [31:0] io_data_writeAddr_bits_addr,
  output [3:0]  io_data_writeAddr_bits_id,
  output [2:0]  io_data_writeAddr_bits_size,
  output [7:0]  io_data_writeAddr_bits_len,
  output [1:0]  io_data_writeAddr_bits_burst,
  output        io_data_writeAddr_bits_lock,
  output [3:0]  io_data_writeAddr_bits_cache,
  output [2:0]  io_data_writeAddr_bits_prot,
  input         io_data_writeData_ready,
  output        io_data_writeData_valid,
  output [31:0] io_data_writeData_bits_data,
  output [3:0]  io_data_writeData_bits_id,
  output        io_data_writeData_bits_last,
  output [3:0]  io_data_writeData_bits_strb,
  output        io_data_writeResp_ready,
  input         io_data_writeResp_valid,
  input  [3:0]  io_data_writeResp_bits_id,
  input  [1:0]  io_data_writeResp_bits_resp,
  input         io_uncached_readAddr_ready,
  output        io_uncached_readAddr_valid,
  output [31:0] io_uncached_readAddr_bits_addr,
  output [3:0]  io_uncached_readAddr_bits_id,
  output [2:0]  io_uncached_readAddr_bits_size,
  output [7:0]  io_uncached_readAddr_bits_len,
  output [1:0]  io_uncached_readAddr_bits_burst,
  output        io_uncached_readAddr_bits_lock,
  output [3:0]  io_uncached_readAddr_bits_cache,
  output [2:0]  io_uncached_readAddr_bits_prot,
  output        io_uncached_readData_ready,
  input         io_uncached_readData_valid,
  input  [31:0] io_uncached_readData_bits_data,
  input  [3:0]  io_uncached_readData_bits_id,
  input         io_uncached_readData_bits_last,
  input  [1:0]  io_uncached_readData_bits_resp,
  input         io_uncached_writeAddr_ready,
  output        io_uncached_writeAddr_valid,
  output [31:0] io_uncached_writeAddr_bits_addr,
  output [3:0]  io_uncached_writeAddr_bits_id,
  output [2:0]  io_uncached_writeAddr_bits_size,
  output [7:0]  io_uncached_writeAddr_bits_len,
  output [1:0]  io_uncached_writeAddr_bits_burst,
  output        io_uncached_writeAddr_bits_lock,
  output [3:0]  io_uncached_writeAddr_bits_cache,
  output [2:0]  io_uncached_writeAddr_bits_prot,
  input         io_uncached_writeData_ready,
  output        io_uncached_writeData_valid,
  output [31:0] io_uncached_writeData_bits_data,
  output [3:0]  io_uncached_writeData_bits_id,
  output        io_uncached_writeData_bits_last,
  output [3:0]  io_uncached_writeData_bits_strb,
  output        io_uncached_writeResp_ready,
  input         io_uncached_writeResp_valid,
  input  [3:0]  io_uncached_writeResp_bits_id,
  input  [1:0]  io_uncached_writeResp_bits_resp
);
  wire  core_clock; // @[Fuxi.scala 22:23]
  wire  core_reset; // @[Fuxi.scala 22:23]
  wire  core_io_irq_timer; // @[Fuxi.scala 22:23]
  wire  core_io_irq_soft; // @[Fuxi.scala 22:23]
  wire  core_io_irq_extern; // @[Fuxi.scala 22:23]
  wire  core_io_tlb_en; // @[Fuxi.scala 22:23]
  wire  core_io_tlb_flushInst; // @[Fuxi.scala 22:23]
  wire  core_io_tlb_flushData; // @[Fuxi.scala 22:23]
  wire [21:0] core_io_tlb_basePpn; // @[Fuxi.scala 22:23]
  wire  core_io_tlb_sum; // @[Fuxi.scala 22:23]
  wire  core_io_tlb_smode; // @[Fuxi.scala 22:23]
  wire  core_io_cache_flushInst; // @[Fuxi.scala 22:23]
  wire  core_io_cache_flushData; // @[Fuxi.scala 22:23]
  wire  core_io_rom_valid; // @[Fuxi.scala 22:23]
  wire  core_io_rom_fault; // @[Fuxi.scala 22:23]
  wire [31:0] core_io_rom_addr; // @[Fuxi.scala 22:23]
  wire [31:0] core_io_rom_rdata; // @[Fuxi.scala 22:23]
  wire  core_io_ram_en; // @[Fuxi.scala 22:23]
  wire  core_io_ram_valid; // @[Fuxi.scala 22:23]
  wire  core_io_ram_fault; // @[Fuxi.scala 22:23]
  wire [3:0] core_io_ram_wen; // @[Fuxi.scala 22:23]
  wire [31:0] core_io_ram_addr; // @[Fuxi.scala 22:23]
  wire [31:0] core_io_ram_rdata; // @[Fuxi.scala 22:23]
  wire [31:0] core_io_ram_wdata; // @[Fuxi.scala 22:23]
  wire  core_io_debug_regWen; // @[Fuxi.scala 22:23]
  wire [4:0] core_io_debug_regWaddr; // @[Fuxi.scala 22:23]
  wire [31:0] core_io_debug_regWdata; // @[Fuxi.scala 22:23]
  wire [31:0] core_io_debug_pc; // @[Fuxi.scala 22:23]
  wire  coreBus_clock; // @[Fuxi.scala 23:23]
  wire  coreBus_reset; // @[Fuxi.scala 23:23]
  wire  coreBus_io_rom_valid; // @[Fuxi.scala 23:23]
  wire  coreBus_io_rom_fault; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_rom_addr; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_rom_rdata; // @[Fuxi.scala 23:23]
  wire  coreBus_io_ram_en; // @[Fuxi.scala 23:23]
  wire  coreBus_io_ram_valid; // @[Fuxi.scala 23:23]
  wire  coreBus_io_ram_fault; // @[Fuxi.scala 23:23]
  wire [3:0] coreBus_io_ram_wen; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_ram_addr; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_ram_rdata; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_ram_wdata; // @[Fuxi.scala 23:23]
  wire  coreBus_io_tlb_en; // @[Fuxi.scala 23:23]
  wire  coreBus_io_tlb_flushInst; // @[Fuxi.scala 23:23]
  wire  coreBus_io_tlb_flushData; // @[Fuxi.scala 23:23]
  wire [21:0] coreBus_io_tlb_basePpn; // @[Fuxi.scala 23:23]
  wire  coreBus_io_tlb_sum; // @[Fuxi.scala 23:23]
  wire  coreBus_io_tlb_smode; // @[Fuxi.scala 23:23]
  wire  coreBus_io_cache_flushInst; // @[Fuxi.scala 23:23]
  wire  coreBus_io_cache_flushData; // @[Fuxi.scala 23:23]
  wire  coreBus_io_inst_readAddr_ready; // @[Fuxi.scala 23:23]
  wire  coreBus_io_inst_readAddr_valid; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_inst_readAddr_bits_addr; // @[Fuxi.scala 23:23]
  wire  coreBus_io_inst_readData_valid; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_inst_readData_bits_data; // @[Fuxi.scala 23:23]
  wire  coreBus_io_inst_readData_bits_last; // @[Fuxi.scala 23:23]
  wire  coreBus_io_data_readAddr_ready; // @[Fuxi.scala 23:23]
  wire  coreBus_io_data_readAddr_valid; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_data_readAddr_bits_addr; // @[Fuxi.scala 23:23]
  wire  coreBus_io_data_readData_valid; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_data_readData_bits_data; // @[Fuxi.scala 23:23]
  wire  coreBus_io_data_readData_bits_last; // @[Fuxi.scala 23:23]
  wire  coreBus_io_data_writeAddr_ready; // @[Fuxi.scala 23:23]
  wire  coreBus_io_data_writeAddr_valid; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_data_writeAddr_bits_addr; // @[Fuxi.scala 23:23]
  wire  coreBus_io_data_writeData_ready; // @[Fuxi.scala 23:23]
  wire  coreBus_io_data_writeData_valid; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_data_writeData_bits_data; // @[Fuxi.scala 23:23]
  wire  coreBus_io_data_writeData_bits_last; // @[Fuxi.scala 23:23]
  wire  coreBus_io_uncached_readAddr_ready; // @[Fuxi.scala 23:23]
  wire  coreBus_io_uncached_readAddr_valid; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_uncached_readAddr_bits_addr; // @[Fuxi.scala 23:23]
  wire  coreBus_io_uncached_readData_valid; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_uncached_readData_bits_data; // @[Fuxi.scala 23:23]
  wire  coreBus_io_uncached_readData_bits_last; // @[Fuxi.scala 23:23]
  wire  coreBus_io_uncached_writeAddr_ready; // @[Fuxi.scala 23:23]
  wire  coreBus_io_uncached_writeAddr_valid; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_uncached_writeAddr_bits_addr; // @[Fuxi.scala 23:23]
  wire  coreBus_io_uncached_writeData_ready; // @[Fuxi.scala 23:23]
  wire  coreBus_io_uncached_writeData_valid; // @[Fuxi.scala 23:23]
  wire [31:0] coreBus_io_uncached_writeData_bits_data; // @[Fuxi.scala 23:23]
  wire  coreBus_io_uncached_writeData_bits_last; // @[Fuxi.scala 23:23]
  wire [3:0] coreBus_io_uncached_writeData_bits_strb; // @[Fuxi.scala 23:23]
  Core core ( // @[Fuxi.scala 22:23]
    .clock(core_clock),
    .reset(core_reset),
    .io_irq_timer(core_io_irq_timer),
    .io_irq_soft(core_io_irq_soft),
    .io_irq_extern(core_io_irq_extern),
    .io_tlb_en(core_io_tlb_en),
    .io_tlb_flushInst(core_io_tlb_flushInst),
    .io_tlb_flushData(core_io_tlb_flushData),
    .io_tlb_basePpn(core_io_tlb_basePpn),
    .io_tlb_sum(core_io_tlb_sum),
    .io_tlb_smode(core_io_tlb_smode),
    .io_cache_flushInst(core_io_cache_flushInst),
    .io_cache_flushData(core_io_cache_flushData),
    .io_rom_valid(core_io_rom_valid),
    .io_rom_fault(core_io_rom_fault),
    .io_rom_addr(core_io_rom_addr),
    .io_rom_rdata(core_io_rom_rdata),
    .io_ram_en(core_io_ram_en),
    .io_ram_valid(core_io_ram_valid),
    .io_ram_fault(core_io_ram_fault),
    .io_ram_wen(core_io_ram_wen),
    .io_ram_addr(core_io_ram_addr),
    .io_ram_rdata(core_io_ram_rdata),
    .io_ram_wdata(core_io_ram_wdata),
    .io_debug_regWen(core_io_debug_regWen),
    .io_debug_regWaddr(core_io_debug_regWaddr),
    .io_debug_regWdata(core_io_debug_regWdata),
    .io_debug_pc(core_io_debug_pc)
  );
  CoreBus coreBus ( // @[Fuxi.scala 23:23]
    .clock(coreBus_clock),
    .reset(coreBus_reset),
    .io_rom_valid(coreBus_io_rom_valid),
    .io_rom_fault(coreBus_io_rom_fault),
    .io_rom_addr(coreBus_io_rom_addr),
    .io_rom_rdata(coreBus_io_rom_rdata),
    .io_ram_en(coreBus_io_ram_en),
    .io_ram_valid(coreBus_io_ram_valid),
    .io_ram_fault(coreBus_io_ram_fault),
    .io_ram_wen(coreBus_io_ram_wen),
    .io_ram_addr(coreBus_io_ram_addr),
    .io_ram_rdata(coreBus_io_ram_rdata),
    .io_ram_wdata(coreBus_io_ram_wdata),
    .io_tlb_en(coreBus_io_tlb_en),
    .io_tlb_flushInst(coreBus_io_tlb_flushInst),
    .io_tlb_flushData(coreBus_io_tlb_flushData),
    .io_tlb_basePpn(coreBus_io_tlb_basePpn),
    .io_tlb_sum(coreBus_io_tlb_sum),
    .io_tlb_smode(coreBus_io_tlb_smode),
    .io_cache_flushInst(coreBus_io_cache_flushInst),
    .io_cache_flushData(coreBus_io_cache_flushData),
    .io_inst_readAddr_ready(coreBus_io_inst_readAddr_ready),
    .io_inst_readAddr_valid(coreBus_io_inst_readAddr_valid),
    .io_inst_readAddr_bits_addr(coreBus_io_inst_readAddr_bits_addr),
    .io_inst_readData_valid(coreBus_io_inst_readData_valid),
    .io_inst_readData_bits_data(coreBus_io_inst_readData_bits_data),
    .io_inst_readData_bits_last(coreBus_io_inst_readData_bits_last),
    .io_data_readAddr_ready(coreBus_io_data_readAddr_ready),
    .io_data_readAddr_valid(coreBus_io_data_readAddr_valid),
    .io_data_readAddr_bits_addr(coreBus_io_data_readAddr_bits_addr),
    .io_data_readData_valid(coreBus_io_data_readData_valid),
    .io_data_readData_bits_data(coreBus_io_data_readData_bits_data),
    .io_data_readData_bits_last(coreBus_io_data_readData_bits_last),
    .io_data_writeAddr_ready(coreBus_io_data_writeAddr_ready),
    .io_data_writeAddr_valid(coreBus_io_data_writeAddr_valid),
    .io_data_writeAddr_bits_addr(coreBus_io_data_writeAddr_bits_addr),
    .io_data_writeData_ready(coreBus_io_data_writeData_ready),
    .io_data_writeData_valid(coreBus_io_data_writeData_valid),
    .io_data_writeData_bits_data(coreBus_io_data_writeData_bits_data),
    .io_data_writeData_bits_last(coreBus_io_data_writeData_bits_last),
    .io_uncached_readAddr_ready(coreBus_io_uncached_readAddr_ready),
    .io_uncached_readAddr_valid(coreBus_io_uncached_readAddr_valid),
    .io_uncached_readAddr_bits_addr(coreBus_io_uncached_readAddr_bits_addr),
    .io_uncached_readData_valid(coreBus_io_uncached_readData_valid),
    .io_uncached_readData_bits_data(coreBus_io_uncached_readData_bits_data),
    .io_uncached_readData_bits_last(coreBus_io_uncached_readData_bits_last),
    .io_uncached_writeAddr_ready(coreBus_io_uncached_writeAddr_ready),
    .io_uncached_writeAddr_valid(coreBus_io_uncached_writeAddr_valid),
    .io_uncached_writeAddr_bits_addr(coreBus_io_uncached_writeAddr_bits_addr),
    .io_uncached_writeData_ready(coreBus_io_uncached_writeData_ready),
    .io_uncached_writeData_valid(coreBus_io_uncached_writeData_valid),
    .io_uncached_writeData_bits_data(coreBus_io_uncached_writeData_bits_data),
    .io_uncached_writeData_bits_last(coreBus_io_uncached_writeData_bits_last),
    .io_uncached_writeData_bits_strb(coreBus_io_uncached_writeData_bits_strb)
  );
  assign io_debug_regWen = core_io_debug_regWen; // @[Fuxi.scala 30:17]
  assign io_debug_regWaddr = core_io_debug_regWaddr; // @[Fuxi.scala 30:17]
  assign io_debug_regWdata = core_io_debug_regWdata; // @[Fuxi.scala 30:17]
  assign io_debug_pc = core_io_debug_pc; // @[Fuxi.scala 30:17]
  assign io_inst_readAddr_valid = coreBus_io_inst_readAddr_valid; // @[Fuxi.scala 32:23]
  assign io_inst_readAddr_bits_addr = coreBus_io_inst_readAddr_bits_addr; // @[Fuxi.scala 32:23]
  assign io_inst_readAddr_bits_id = 4'h0; // @[Fuxi.scala 32:23]
  assign io_inst_readAddr_bits_size = 3'h2; // @[Fuxi.scala 32:23]
  assign io_inst_readAddr_bits_len = 8'hf; // @[Fuxi.scala 32:23]
  assign io_inst_readAddr_bits_burst = 2'h1; // @[Fuxi.scala 32:23]
  assign io_inst_readAddr_bits_lock = 1'h0; // @[Fuxi.scala 32:23]
  assign io_inst_readAddr_bits_cache = 4'h0; // @[Fuxi.scala 32:23]
  assign io_inst_readAddr_bits_prot = 3'h0; // @[Fuxi.scala 32:23]
  assign io_inst_readData_ready = 1'h1; // @[Fuxi.scala 32:23]
  assign io_inst_writeAddr_valid = 1'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeAddr_bits_addr = 32'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeAddr_bits_id = 4'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeAddr_bits_size = 3'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeAddr_bits_len = 8'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeAddr_bits_burst = 2'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeAddr_bits_lock = 1'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeAddr_bits_cache = 4'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeAddr_bits_prot = 3'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeData_valid = 1'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeData_bits_data = 32'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeData_bits_id = 4'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeData_bits_last = 1'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeData_bits_strb = 4'h0; // @[Fuxi.scala 32:23]
  assign io_inst_writeResp_ready = 1'h0; // @[Fuxi.scala 32:23]
  assign io_data_readAddr_valid = coreBus_io_data_readAddr_valid; // @[Fuxi.scala 33:23]
  assign io_data_readAddr_bits_addr = coreBus_io_data_readAddr_bits_addr; // @[Fuxi.scala 33:23]
  assign io_data_readAddr_bits_id = 4'h0; // @[Fuxi.scala 33:23]
  assign io_data_readAddr_bits_size = 3'h2; // @[Fuxi.scala 33:23]
  assign io_data_readAddr_bits_len = 8'hf; // @[Fuxi.scala 33:23]
  assign io_data_readAddr_bits_burst = 2'h1; // @[Fuxi.scala 33:23]
  assign io_data_readAddr_bits_lock = 1'h0; // @[Fuxi.scala 33:23]
  assign io_data_readAddr_bits_cache = 4'h0; // @[Fuxi.scala 33:23]
  assign io_data_readAddr_bits_prot = 3'h0; // @[Fuxi.scala 33:23]
  assign io_data_readData_ready = 1'h1; // @[Fuxi.scala 33:23]
  assign io_data_writeAddr_valid = coreBus_io_data_writeAddr_valid; // @[Fuxi.scala 33:23]
  assign io_data_writeAddr_bits_addr = coreBus_io_data_writeAddr_bits_addr; // @[Fuxi.scala 33:23]
  assign io_data_writeAddr_bits_id = 4'h0; // @[Fuxi.scala 33:23]
  assign io_data_writeAddr_bits_size = 3'h2; // @[Fuxi.scala 33:23]
  assign io_data_writeAddr_bits_len = 8'hf; // @[Fuxi.scala 33:23]
  assign io_data_writeAddr_bits_burst = 2'h1; // @[Fuxi.scala 33:23]
  assign io_data_writeAddr_bits_lock = 1'h0; // @[Fuxi.scala 33:23]
  assign io_data_writeAddr_bits_cache = 4'h0; // @[Fuxi.scala 33:23]
  assign io_data_writeAddr_bits_prot = 3'h0; // @[Fuxi.scala 33:23]
  assign io_data_writeData_valid = coreBus_io_data_writeData_valid; // @[Fuxi.scala 33:23]
  assign io_data_writeData_bits_data = coreBus_io_data_writeData_bits_data; // @[Fuxi.scala 33:23]
  assign io_data_writeData_bits_id = 4'h0; // @[Fuxi.scala 33:23]
  assign io_data_writeData_bits_last = coreBus_io_data_writeData_bits_last; // @[Fuxi.scala 33:23]
  assign io_data_writeData_bits_strb = 4'hf; // @[Fuxi.scala 33:23]
  assign io_data_writeResp_ready = 1'h1; // @[Fuxi.scala 33:23]
  assign io_uncached_readAddr_valid = coreBus_io_uncached_readAddr_valid; // @[Fuxi.scala 34:23]
  assign io_uncached_readAddr_bits_addr = coreBus_io_uncached_readAddr_bits_addr; // @[Fuxi.scala 34:23]
  assign io_uncached_readAddr_bits_id = 4'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_readAddr_bits_size = 3'h2; // @[Fuxi.scala 34:23]
  assign io_uncached_readAddr_bits_len = 8'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_readAddr_bits_burst = 2'h1; // @[Fuxi.scala 34:23]
  assign io_uncached_readAddr_bits_lock = 1'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_readAddr_bits_cache = 4'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_readAddr_bits_prot = 3'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_readData_ready = 1'h1; // @[Fuxi.scala 34:23]
  assign io_uncached_writeAddr_valid = coreBus_io_uncached_writeAddr_valid; // @[Fuxi.scala 34:23]
  assign io_uncached_writeAddr_bits_addr = coreBus_io_uncached_writeAddr_bits_addr; // @[Fuxi.scala 34:23]
  assign io_uncached_writeAddr_bits_id = 4'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_writeAddr_bits_size = 3'h2; // @[Fuxi.scala 34:23]
  assign io_uncached_writeAddr_bits_len = 8'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_writeAddr_bits_burst = 2'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_writeAddr_bits_lock = 1'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_writeAddr_bits_cache = 4'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_writeAddr_bits_prot = 3'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_writeData_valid = coreBus_io_uncached_writeData_valid; // @[Fuxi.scala 34:23]
  assign io_uncached_writeData_bits_data = coreBus_io_uncached_writeData_bits_data; // @[Fuxi.scala 34:23]
  assign io_uncached_writeData_bits_id = 4'h0; // @[Fuxi.scala 34:23]
  assign io_uncached_writeData_bits_last = coreBus_io_uncached_writeData_bits_last; // @[Fuxi.scala 34:23]
  assign io_uncached_writeData_bits_strb = coreBus_io_uncached_writeData_bits_strb; // @[Fuxi.scala 34:23]
  assign io_uncached_writeResp_ready = 1'h1; // @[Fuxi.scala 34:23]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_irq_timer = io_irq_timer; // @[Fuxi.scala 25:17]
  assign core_io_irq_soft = io_irq_soft; // @[Fuxi.scala 25:17]
  assign core_io_irq_extern = io_irq_extern; // @[Fuxi.scala 25:17]
  assign core_io_rom_valid = coreBus_io_rom_valid; // @[Fuxi.scala 28:17]
  assign core_io_rom_fault = coreBus_io_rom_fault; // @[Fuxi.scala 28:17]
  assign core_io_rom_rdata = coreBus_io_rom_rdata; // @[Fuxi.scala 28:17]
  assign core_io_ram_valid = coreBus_io_ram_valid; // @[Fuxi.scala 29:17]
  assign core_io_ram_fault = coreBus_io_ram_fault; // @[Fuxi.scala 29:17]
  assign core_io_ram_rdata = coreBus_io_ram_rdata; // @[Fuxi.scala 29:17]
  assign coreBus_clock = clock;
  assign coreBus_reset = reset;
  assign coreBus_io_rom_addr = core_io_rom_addr; // @[Fuxi.scala 28:17]
  assign coreBus_io_ram_en = core_io_ram_en; // @[Fuxi.scala 29:17]
  assign coreBus_io_ram_wen = core_io_ram_wen; // @[Fuxi.scala 29:17]
  assign coreBus_io_ram_addr = core_io_ram_addr; // @[Fuxi.scala 29:17]
  assign coreBus_io_ram_wdata = core_io_ram_wdata; // @[Fuxi.scala 29:17]
  assign coreBus_io_tlb_en = core_io_tlb_en; // @[Fuxi.scala 26:17]
  assign coreBus_io_tlb_flushInst = core_io_tlb_flushInst; // @[Fuxi.scala 26:17]
  assign coreBus_io_tlb_flushData = core_io_tlb_flushData; // @[Fuxi.scala 26:17]
  assign coreBus_io_tlb_basePpn = core_io_tlb_basePpn; // @[Fuxi.scala 26:17]
  assign coreBus_io_tlb_sum = core_io_tlb_sum; // @[Fuxi.scala 26:17]
  assign coreBus_io_tlb_smode = core_io_tlb_smode; // @[Fuxi.scala 26:17]
  assign coreBus_io_cache_flushInst = core_io_cache_flushInst; // @[Fuxi.scala 27:17]
  assign coreBus_io_cache_flushData = core_io_cache_flushData; // @[Fuxi.scala 27:17]
  assign coreBus_io_inst_readAddr_ready = io_inst_readAddr_ready; // @[Fuxi.scala 32:23]
  assign coreBus_io_inst_readData_valid = io_inst_readData_valid; // @[Fuxi.scala 32:23]
  assign coreBus_io_inst_readData_bits_data = io_inst_readData_bits_data; // @[Fuxi.scala 32:23]
  assign coreBus_io_inst_readData_bits_last = io_inst_readData_bits_last; // @[Fuxi.scala 32:23]
  assign coreBus_io_data_readAddr_ready = io_data_readAddr_ready; // @[Fuxi.scala 33:23]
  assign coreBus_io_data_readData_valid = io_data_readData_valid; // @[Fuxi.scala 33:23]
  assign coreBus_io_data_readData_bits_data = io_data_readData_bits_data; // @[Fuxi.scala 33:23]
  assign coreBus_io_data_readData_bits_last = io_data_readData_bits_last; // @[Fuxi.scala 33:23]
  assign coreBus_io_data_writeAddr_ready = io_data_writeAddr_ready; // @[Fuxi.scala 33:23]
  assign coreBus_io_data_writeData_ready = io_data_writeData_ready; // @[Fuxi.scala 33:23]
  assign coreBus_io_uncached_readAddr_ready = io_uncached_readAddr_ready; // @[Fuxi.scala 34:23]
  assign coreBus_io_uncached_readData_valid = io_uncached_readData_valid; // @[Fuxi.scala 34:23]
  assign coreBus_io_uncached_readData_bits_data = io_uncached_readData_bits_data; // @[Fuxi.scala 34:23]
  assign coreBus_io_uncached_readData_bits_last = io_uncached_readData_bits_last; // @[Fuxi.scala 34:23]
  assign coreBus_io_uncached_writeAddr_ready = io_uncached_writeAddr_ready; // @[Fuxi.scala 34:23]
  assign coreBus_io_uncached_writeData_ready = io_uncached_writeData_ready; // @[Fuxi.scala 34:23]
endmodule
